module CSRFile( // @[:@2591.2]
  input         clock, // @[:@2592.4]
  input         reset, // @[:@2593.4]
  input  [2:0]  io_rw_cmd, // @[:@2594.4]
  input  [11:0] io_rw_addr, // @[:@2594.4]
  output [31:0] io_rw_rdata, // @[:@2594.4]
  input  [31:0] io_rw_wdata, // @[:@2594.4]
  output        io_eret, // @[:@2594.4]
  output [1:0]  io_status_prv, // @[:@2594.4]
  output [13:0] io_status_unimp5, // @[:@2594.4]
  output        io_status_mprv, // @[:@2594.4]
  output [1:0]  io_status_unimp4, // @[:@2594.4]
  output [1:0]  io_status_mpp, // @[:@2594.4]
  output [2:0]  io_status_unimp3, // @[:@2594.4]
  output        io_status_mpie, // @[:@2594.4]
  output [2:0]  io_status_unimp2, // @[:@2594.4]
  output        io_status_mie, // @[:@2594.4]
  output [2:0]  io_status_unimp1, // @[:@2594.4]
  input         io_xcpt, // @[:@2594.4]
  input  [31:0] io_cause, // @[:@2594.4]
  input  [31:0] io_tval, // @[:@2594.4]
  output [31:0] io_evec, // @[:@2594.4]
  input         io_illegal, // @[:@2594.4]
  input  [1:0]  io_retire, // @[:@2594.4]
  input  [31:0] io_pc, // @[:@2594.4]
  output [31:0] io_time // @[:@2594.4]
);
  reg [1:0] reg_mstatus_prv; // @[CSR.scala 112:28:@2721.4]
  reg [31:0] _RAND_0;
  reg  reg_mstatus_mpie; // @[CSR.scala 112:28:@2721.4]
  reg [31:0] _RAND_1;
  reg  reg_mstatus_mie; // @[CSR.scala 112:28:@2721.4]
  reg [31:0] _RAND_2;
  reg [31:0] reg_mepc; // @[CSR.scala 113:21:@2722.4]
  reg [31:0] _RAND_3;
  reg [31:0] reg_mcause; // @[CSR.scala 114:23:@2723.4]
  reg [31:0] _RAND_4;
  reg [31:0] reg_mtval; // @[CSR.scala 115:22:@2724.4]
  reg [31:0] _RAND_5;
  reg [31:0] reg_mscratch; // @[CSR.scala 116:25:@2725.4]
  reg [31:0] _RAND_6;
  reg [31:0] reg_medeleg; // @[CSR.scala 118:24:@2727.4]
  reg [31:0] _RAND_7;
  reg  reg_mip_mtip; // @[CSR.scala 120:24:@2745.4]
  reg [31:0] _RAND_8;
  reg  reg_mip_msip; // @[CSR.scala 120:24:@2745.4]
  reg [31:0] _RAND_9;
  reg  reg_mie_mtip; // @[CSR.scala 121:24:@2763.4]
  reg [31:0] _RAND_10;
  reg  reg_mie_msip; // @[CSR.scala 121:24:@2763.4]
  reg [31:0] _RAND_11;
  reg [5:0] _T_240; // @[Util.scala 112:41:@2766.4]
  reg [31:0] _RAND_12;
  wire [6:0] _T_241; // @[Util.scala 113:33:@2767.4]
  reg [57:0] _T_244; // @[Util.scala 117:31:@2769.4]
  reg [63:0] _RAND_13;
  wire  _T_245; // @[Util.scala 118:20:@2770.4]
  wire [58:0] _T_247; // @[Util.scala 118:43:@2772.6]
  wire [57:0] _T_248; // @[Util.scala 118:43:@2773.6]
  wire [57:0] _GEN_0; // @[Util.scala 118:34:@2771.4]
  wire [63:0] _T_249; // @[Cat.scala 30:58:@2776.4]
  reg [5:0] _T_252; // @[Util.scala 112:41:@2777.4]
  reg [31:0] _RAND_14;
  wire [5:0] _GEN_147; // @[Util.scala 113:33:@2778.4]
  wire [6:0] _T_253; // @[Util.scala 113:33:@2778.4]
  reg [57:0] _T_256; // @[Util.scala 117:31:@2780.4]
  reg [63:0] _RAND_15;
  wire  _T_257; // @[Util.scala 118:20:@2781.4]
  wire [58:0] _T_259; // @[Util.scala 118:43:@2783.6]
  wire [57:0] _T_260; // @[Util.scala 118:43:@2784.6]
  wire [57:0] _GEN_1; // @[Util.scala 118:34:@2782.4]
  wire [63:0] _T_261; // @[Cat.scala 30:58:@2787.4]
  reg [39:0] _T_264; // @[Util.scala 112:74:@2789.4]
  reg [63:0] _RAND_16;
  wire [40:0] _T_265; // @[Util.scala 113:33:@2790.4]
  reg [39:0] _T_267; // @[Util.scala 112:74:@2792.4]
  reg [63:0] _RAND_17;
  wire [40:0] _T_268; // @[Util.scala 113:33:@2793.4]
  reg [39:0] _T_270; // @[Util.scala 112:74:@2795.4]
  reg [63:0] _RAND_18;
  wire [40:0] _T_271; // @[Util.scala 113:33:@2796.4]
  reg [39:0] _T_273; // @[Util.scala 112:74:@2798.4]
  reg [63:0] _RAND_19;
  wire [40:0] _T_274; // @[Util.scala 113:33:@2799.4]
  reg [39:0] _T_276; // @[Util.scala 112:74:@2801.4]
  reg [63:0] _RAND_20;
  wire [40:0] _T_277; // @[Util.scala 113:33:@2802.4]
  reg [39:0] _T_279; // @[Util.scala 112:74:@2804.4]
  reg [63:0] _RAND_21;
  wire [40:0] _T_280; // @[Util.scala 113:33:@2805.4]
  reg [39:0] _T_282; // @[Util.scala 112:74:@2807.4]
  reg [63:0] _RAND_22;
  wire [40:0] _T_283; // @[Util.scala 113:33:@2808.4]
  reg [39:0] _T_285; // @[Util.scala 112:74:@2810.4]
  reg [63:0] _RAND_23;
  wire [40:0] _T_286; // @[Util.scala 113:33:@2811.4]
  reg [39:0] _T_288; // @[Util.scala 112:74:@2813.4]
  reg [63:0] _RAND_24;
  wire [40:0] _T_289; // @[Util.scala 113:33:@2814.4]
  reg [39:0] _T_291; // @[Util.scala 112:74:@2816.4]
  reg [63:0] _RAND_25;
  wire [40:0] _T_292; // @[Util.scala 113:33:@2817.4]
  reg [39:0] _T_294; // @[Util.scala 112:74:@2819.4]
  reg [63:0] _RAND_26;
  wire [40:0] _T_295; // @[Util.scala 113:33:@2820.4]
  reg [39:0] _T_297; // @[Util.scala 112:74:@2822.4]
  reg [63:0] _RAND_27;
  wire [40:0] _T_298; // @[Util.scala 113:33:@2823.4]
  reg [39:0] _T_300; // @[Util.scala 112:74:@2825.4]
  reg [63:0] _RAND_28;
  wire [40:0] _T_301; // @[Util.scala 113:33:@2826.4]
  reg [39:0] _T_303; // @[Util.scala 112:74:@2828.4]
  reg [63:0] _RAND_29;
  wire [40:0] _T_304; // @[Util.scala 113:33:@2829.4]
  reg [39:0] _T_306; // @[Util.scala 112:74:@2831.4]
  reg [63:0] _RAND_30;
  wire [40:0] _T_307; // @[Util.scala 113:33:@2832.4]
  reg [39:0] _T_309; // @[Util.scala 112:74:@2834.4]
  reg [63:0] _RAND_31;
  wire [40:0] _T_310; // @[Util.scala 113:33:@2835.4]
  reg [39:0] _T_312; // @[Util.scala 112:74:@2837.4]
  reg [63:0] _RAND_32;
  wire [40:0] _T_313; // @[Util.scala 113:33:@2838.4]
  reg [39:0] _T_315; // @[Util.scala 112:74:@2840.4]
  reg [63:0] _RAND_33;
  wire [40:0] _T_316; // @[Util.scala 113:33:@2841.4]
  reg [39:0] _T_318; // @[Util.scala 112:74:@2843.4]
  reg [63:0] _RAND_34;
  wire [40:0] _T_319; // @[Util.scala 113:33:@2844.4]
  reg [39:0] _T_321; // @[Util.scala 112:74:@2846.4]
  reg [63:0] _RAND_35;
  wire [40:0] _T_322; // @[Util.scala 113:33:@2847.4]
  reg [39:0] _T_324; // @[Util.scala 112:74:@2849.4]
  reg [63:0] _RAND_36;
  wire [40:0] _T_325; // @[Util.scala 113:33:@2850.4]
  reg [39:0] _T_327; // @[Util.scala 112:74:@2852.4]
  reg [63:0] _RAND_37;
  wire [40:0] _T_328; // @[Util.scala 113:33:@2853.4]
  reg [39:0] _T_330; // @[Util.scala 112:74:@2855.4]
  reg [63:0] _RAND_38;
  wire [40:0] _T_331; // @[Util.scala 113:33:@2856.4]
  reg [39:0] _T_333; // @[Util.scala 112:74:@2858.4]
  reg [63:0] _RAND_39;
  wire [40:0] _T_334; // @[Util.scala 113:33:@2859.4]
  reg [39:0] _T_336; // @[Util.scala 112:74:@2861.4]
  reg [63:0] _RAND_40;
  wire [40:0] _T_337; // @[Util.scala 113:33:@2862.4]
  reg [39:0] _T_339; // @[Util.scala 112:74:@2864.4]
  reg [63:0] _RAND_41;
  wire [40:0] _T_340; // @[Util.scala 113:33:@2865.4]
  reg [39:0] _T_342; // @[Util.scala 112:74:@2867.4]
  reg [63:0] _RAND_42;
  wire [40:0] _T_343; // @[Util.scala 113:33:@2868.4]
  reg [39:0] _T_345; // @[Util.scala 112:74:@2870.4]
  reg [63:0] _RAND_43;
  wire [40:0] _T_346; // @[Util.scala 113:33:@2871.4]
  reg [39:0] _T_348; // @[Util.scala 112:74:@2873.4]
  reg [63:0] _RAND_44;
  wire [40:0] _T_349; // @[Util.scala 113:33:@2874.4]
  reg [39:0] _T_351; // @[Util.scala 112:74:@2876.4]
  reg [63:0] _RAND_45;
  wire [40:0] _T_352; // @[Util.scala 113:33:@2877.4]
  reg [39:0] _T_354; // @[Util.scala 112:74:@2879.4]
  reg [63:0] _RAND_46;
  wire [40:0] _T_355; // @[Util.scala 113:33:@2880.4]
  reg [39:0] _T_357; // @[Util.scala 112:74:@2882.4]
  reg [63:0] _RAND_47;
  wire [40:0] _T_358; // @[Util.scala 113:33:@2883.4]
  reg [31:0] reg_dscratch; // @[CSR.scala 134:25:@2972.4]
  reg [31:0] _RAND_48;
  wire  system_insn; // @[CSR.scala 137:31:@2974.4]
  wire  _T_446; // @[CSR.scala 138:27:@2975.4]
  wire  _T_448; // @[CSR.scala 138:40:@2976.4]
  wire  cpu_ren; // @[CSR.scala 138:37:@2977.4]
  wire [31:0] read_mstatus; // @[CSR.scala 140:32:@2986.4]
  wire [15:0] _T_468; // @[CSR.scala 156:25:@2992.4]
  wire [15:0] _T_474; // @[CSR.scala 157:25:@2998.4]
  wire  _T_478; // @[CSR.scala 177:73:@2999.4]
  wire  _T_480; // @[CSR.scala 177:73:@3000.4]
  wire  _T_482; // @[CSR.scala 177:73:@3001.4]
  wire  _T_488; // @[CSR.scala 177:73:@3004.4]
  wire  _T_490; // @[CSR.scala 177:73:@3005.4]
  wire  _T_492; // @[CSR.scala 177:73:@3006.4]
  wire  _T_494; // @[CSR.scala 177:73:@3007.4]
  wire  _T_496; // @[CSR.scala 177:73:@3008.4]
  wire  _T_498; // @[CSR.scala 177:73:@3009.4]
  wire  _T_500; // @[CSR.scala 177:73:@3010.4]
  wire  _T_502; // @[CSR.scala 177:73:@3011.4]
  wire  _T_504; // @[CSR.scala 177:73:@3012.4]
  wire  _T_508; // @[CSR.scala 177:73:@3014.4]
  wire  _T_510; // @[CSR.scala 177:73:@3015.4]
  wire  _T_512; // @[CSR.scala 177:73:@3016.4]
  wire  _T_514; // @[CSR.scala 177:73:@3017.4]
  wire  _T_516; // @[CSR.scala 177:73:@3018.4]
  wire  _T_518; // @[CSR.scala 177:73:@3019.4]
  wire  _T_520; // @[CSR.scala 177:73:@3020.4]
  wire  _T_522; // @[CSR.scala 177:73:@3021.4]
  wire  _T_524; // @[CSR.scala 177:73:@3022.4]
  wire  _T_526; // @[CSR.scala 177:73:@3023.4]
  wire  _T_528; // @[CSR.scala 177:73:@3024.4]
  wire  _T_530; // @[CSR.scala 177:73:@3025.4]
  wire  _T_532; // @[CSR.scala 177:73:@3026.4]
  wire  _T_534; // @[CSR.scala 177:73:@3027.4]
  wire  _T_536; // @[CSR.scala 177:73:@3028.4]
  wire  _T_538; // @[CSR.scala 177:73:@3029.4]
  wire  _T_540; // @[CSR.scala 177:73:@3030.4]
  wire  _T_542; // @[CSR.scala 177:73:@3031.4]
  wire  _T_544; // @[CSR.scala 177:73:@3032.4]
  wire  _T_546; // @[CSR.scala 177:73:@3033.4]
  wire  _T_548; // @[CSR.scala 177:73:@3034.4]
  wire  _T_550; // @[CSR.scala 177:73:@3035.4]
  wire  _T_552; // @[CSR.scala 177:73:@3036.4]
  wire  _T_554; // @[CSR.scala 177:73:@3037.4]
  wire  _T_556; // @[CSR.scala 177:73:@3038.4]
  wire  _T_558; // @[CSR.scala 177:73:@3039.4]
  wire  _T_560; // @[CSR.scala 177:73:@3040.4]
  wire  _T_562; // @[CSR.scala 177:73:@3041.4]
  wire  _T_564; // @[CSR.scala 177:73:@3042.4]
  wire  _T_566; // @[CSR.scala 177:73:@3043.4]
  wire  _T_568; // @[CSR.scala 177:73:@3044.4]
  wire  _T_570; // @[CSR.scala 177:73:@3045.4]
  wire  _T_572; // @[CSR.scala 177:73:@3046.4]
  wire  _T_574; // @[CSR.scala 177:73:@3047.4]
  wire  _T_576; // @[CSR.scala 177:73:@3048.4]
  wire  _T_578; // @[CSR.scala 177:73:@3049.4]
  wire  _T_580; // @[CSR.scala 177:73:@3050.4]
  wire  _T_582; // @[CSR.scala 177:73:@3051.4]
  wire  _T_584; // @[CSR.scala 177:73:@3052.4]
  wire  _T_586; // @[CSR.scala 177:73:@3053.4]
  wire  _T_588; // @[CSR.scala 177:73:@3054.4]
  wire  _T_590; // @[CSR.scala 177:73:@3055.4]
  wire  _T_592; // @[CSR.scala 177:73:@3056.4]
  wire  _T_594; // @[CSR.scala 177:73:@3057.4]
  wire  _T_596; // @[CSR.scala 177:73:@3058.4]
  wire  _T_598; // @[CSR.scala 177:73:@3059.4]
  wire  _T_600; // @[CSR.scala 177:73:@3060.4]
  wire  _T_602; // @[CSR.scala 177:73:@3061.4]
  wire  _T_604; // @[CSR.scala 177:73:@3062.4]
  wire  _T_606; // @[CSR.scala 177:73:@3063.4]
  wire  _T_608; // @[CSR.scala 177:73:@3064.4]
  wire  _T_610; // @[CSR.scala 177:73:@3065.4]
  wire  _T_612; // @[CSR.scala 177:73:@3066.4]
  wire  _T_614; // @[CSR.scala 177:73:@3067.4]
  wire  _T_616; // @[CSR.scala 177:73:@3068.4]
  wire  _T_618; // @[CSR.scala 177:73:@3069.4]
  wire  _T_620; // @[CSR.scala 177:73:@3070.4]
  wire  _T_622; // @[CSR.scala 177:73:@3071.4]
  wire  _T_624; // @[CSR.scala 177:73:@3072.4]
  wire  _T_626; // @[CSR.scala 177:73:@3073.4]
  wire  _T_628; // @[CSR.scala 177:73:@3074.4]
  wire  _T_630; // @[CSR.scala 177:73:@3075.4]
  wire  _T_632; // @[CSR.scala 177:73:@3076.4]
  wire  _T_634; // @[CSR.scala 177:73:@3077.4]
  wire  _T_636; // @[CSR.scala 177:73:@3078.4]
  wire  _T_638; // @[CSR.scala 177:73:@3079.4]
  wire  _T_640; // @[CSR.scala 177:73:@3080.4]
  wire  _T_642; // @[CSR.scala 177:73:@3081.4]
  wire [1:0] _T_643; // @[CSR.scala 179:54:@3082.4]
  wire  priv_sufficient; // @[CSR.scala 179:41:@3083.4]
  wire [1:0] _T_644; // @[CSR.scala 180:29:@3084.4]
  wire [1:0] _T_645; // @[CSR.scala 180:37:@3085.4]
  wire  read_only; // @[CSR.scala 180:37:@3086.4]
  wire  _T_647; // @[CSR.scala 181:38:@3087.4]
  wire  _T_648; // @[CSR.scala 181:25:@3088.4]
  wire  cpu_wen; // @[CSR.scala 181:48:@3089.4]
  wire  _T_650; // @[CSR.scala 182:24:@3090.4]
  wire  wen; // @[CSR.scala 182:21:@3091.4]
  wire  _T_651; // @[Util.scala 23:47:@3092.4]
  wire  _T_652; // @[Util.scala 23:47:@3093.4]
  wire  _T_653; // @[Util.scala 23:62:@3094.4]
  wire [31:0] _T_655; // @[CSR.scala 281:9:@3095.4]
  wire [31:0] _T_656; // @[CSR.scala 281:49:@3096.4]
  wire [31:0] _T_659; // @[CSR.scala 281:64:@3098.4]
  wire [31:0] _T_660; // @[CSR.scala 281:60:@3099.4]
  wire [31:0] wdata; // @[CSR.scala 281:58:@3100.4]
  wire [2:0] _T_662; // @[CSR.scala 185:33:@3101.4]
  wire [7:0] opcode; // @[CSR.scala 185:20:@3102.4]
  wire  _T_663; // @[CSR.scala 186:40:@3103.4]
  wire  insn_call; // @[CSR.scala 186:31:@3104.4]
  wire  _T_664; // @[CSR.scala 187:41:@3105.4]
  wire  insn_break; // @[CSR.scala 187:32:@3106.4]
  wire  _T_665; // @[CSR.scala 188:39:@3107.4]
  wire  _T_666; // @[CSR.scala 188:30:@3108.4]
  wire  insn_ret; // @[CSR.scala 188:43:@3109.4]
  wire  _T_940; // @[CSR.scala 199:24:@3308.4]
  wire [1:0] _T_942; // @[Bitwise.scala 48:55:@3311.4]
  wire  _T_944; // @[CSR.scala 201:50:@3312.4]
  wire  _T_946; // @[CSR.scala 201:9:@3314.4]
  wire  _T_948; // @[CSR.scala 201:9:@3315.4]
  wire  _T_951; // @[CSR.scala 208:32:@3324.4]
  wire  _T_953; // @[CSR.scala 208:21:@3325.4]
  wire  _T_954; // @[CSR.scala 208:18:@3326.4]
  wire  _GEN_3; // @[CSR.scala 208:38:@3327.4]
  wire  _GEN_4; // @[CSR.scala 208:38:@3327.4]
  wire [1:0] new_prv; // @[CSR.scala 208:38:@3327.4]
  wire [3:0] _GEN_148; // @[CSR.scala 218:35:@3335.6]
  wire [4:0] _T_958; // @[CSR.scala 218:35:@3335.6]
  wire [3:0] _T_959; // @[CSR.scala 218:35:@3336.6]
  wire [31:0] _GEN_7; // @[CSR.scala 216:18:@3333.4]
  wire [31:0] _GEN_8; // @[CSR.scala 216:18:@3333.4]
  wire [31:0] _GEN_9; // @[CSR.scala 216:18:@3333.4]
  wire [31:0] _GEN_10; // @[CSR.scala 223:19:@3340.4]
  wire [31:0] _GEN_11; // @[CSR.scala 223:19:@3340.4]
  wire [31:0] _GEN_12; // @[CSR.scala 223:19:@3340.4]
  wire [31:0] _GEN_14; // @[CSR.scala 229:17:@3345.4]
  wire [31:0] _GEN_15; // @[CSR.scala 229:17:@3345.4]
  wire [31:0] _GEN_16; // @[CSR.scala 229:17:@3345.4]
  wire [63:0] _T_965; // @[Mux.scala 19:72:@3353.4]
  wire [63:0] _T_967; // @[Mux.scala 19:72:@3354.4]
  wire [15:0] _T_969; // @[Mux.scala 19:72:@3355.4]
  wire [30:0] _T_975; // @[Mux.scala 19:72:@3358.4]
  wire [31:0] _T_977; // @[Mux.scala 19:72:@3359.4]
  wire [8:0] _T_979; // @[Mux.scala 19:72:@3360.4]
  wire [15:0] _T_981; // @[Mux.scala 19:72:@3361.4]
  wire [15:0] _T_983; // @[Mux.scala 19:72:@3362.4]
  wire [31:0] _T_985; // @[Mux.scala 19:72:@3363.4]
  wire [31:0] _T_987; // @[Mux.scala 19:72:@3364.4]
  wire [31:0] _T_989; // @[Mux.scala 19:72:@3365.4]
  wire [31:0] _T_991; // @[Mux.scala 19:72:@3366.4]
  wire [31:0] _T_995; // @[Mux.scala 19:72:@3368.4]
  wire [31:0] _T_997; // @[Mux.scala 19:72:@3369.4]
  wire [39:0] _T_999; // @[Mux.scala 19:72:@3370.4]
  wire [39:0] _T_1001; // @[Mux.scala 19:72:@3371.4]
  wire [39:0] _T_1003; // @[Mux.scala 19:72:@3372.4]
  wire [39:0] _T_1005; // @[Mux.scala 19:72:@3373.4]
  wire [39:0] _T_1007; // @[Mux.scala 19:72:@3374.4]
  wire [39:0] _T_1009; // @[Mux.scala 19:72:@3375.4]
  wire [39:0] _T_1011; // @[Mux.scala 19:72:@3376.4]
  wire [39:0] _T_1013; // @[Mux.scala 19:72:@3377.4]
  wire [39:0] _T_1015; // @[Mux.scala 19:72:@3378.4]
  wire [39:0] _T_1017; // @[Mux.scala 19:72:@3379.4]
  wire [39:0] _T_1019; // @[Mux.scala 19:72:@3380.4]
  wire [39:0] _T_1021; // @[Mux.scala 19:72:@3381.4]
  wire [39:0] _T_1023; // @[Mux.scala 19:72:@3382.4]
  wire [39:0] _T_1025; // @[Mux.scala 19:72:@3383.4]
  wire [39:0] _T_1027; // @[Mux.scala 19:72:@3384.4]
  wire [39:0] _T_1029; // @[Mux.scala 19:72:@3385.4]
  wire [39:0] _T_1031; // @[Mux.scala 19:72:@3386.4]
  wire [39:0] _T_1033; // @[Mux.scala 19:72:@3387.4]
  wire [39:0] _T_1035; // @[Mux.scala 19:72:@3388.4]
  wire [39:0] _T_1037; // @[Mux.scala 19:72:@3389.4]
  wire [39:0] _T_1039; // @[Mux.scala 19:72:@3390.4]
  wire [39:0] _T_1041; // @[Mux.scala 19:72:@3391.4]
  wire [39:0] _T_1043; // @[Mux.scala 19:72:@3392.4]
  wire [39:0] _T_1045; // @[Mux.scala 19:72:@3393.4]
  wire [39:0] _T_1047; // @[Mux.scala 19:72:@3394.4]
  wire [39:0] _T_1049; // @[Mux.scala 19:72:@3395.4]
  wire [39:0] _T_1051; // @[Mux.scala 19:72:@3396.4]
  wire [39:0] _T_1053; // @[Mux.scala 19:72:@3397.4]
  wire [39:0] _T_1055; // @[Mux.scala 19:72:@3398.4]
  wire [39:0] _T_1057; // @[Mux.scala 19:72:@3399.4]
  wire [39:0] _T_1059; // @[Mux.scala 19:72:@3400.4]
  wire [39:0] _T_1061; // @[Mux.scala 19:72:@3401.4]
  wire [39:0] _T_1063; // @[Mux.scala 19:72:@3402.4]
  wire [39:0] _T_1065; // @[Mux.scala 19:72:@3403.4]
  wire [39:0] _T_1067; // @[Mux.scala 19:72:@3404.4]
  wire [39:0] _T_1069; // @[Mux.scala 19:72:@3405.4]
  wire [39:0] _T_1071; // @[Mux.scala 19:72:@3406.4]
  wire [39:0] _T_1073; // @[Mux.scala 19:72:@3407.4]
  wire [39:0] _T_1075; // @[Mux.scala 19:72:@3408.4]
  wire [39:0] _T_1077; // @[Mux.scala 19:72:@3409.4]
  wire [39:0] _T_1079; // @[Mux.scala 19:72:@3410.4]
  wire [39:0] _T_1081; // @[Mux.scala 19:72:@3411.4]
  wire [39:0] _T_1083; // @[Mux.scala 19:72:@3412.4]
  wire [39:0] _T_1085; // @[Mux.scala 19:72:@3413.4]
  wire [39:0] _T_1087; // @[Mux.scala 19:72:@3414.4]
  wire [39:0] _T_1089; // @[Mux.scala 19:72:@3415.4]
  wire [39:0] _T_1091; // @[Mux.scala 19:72:@3416.4]
  wire [39:0] _T_1093; // @[Mux.scala 19:72:@3417.4]
  wire [39:0] _T_1095; // @[Mux.scala 19:72:@3418.4]
  wire [39:0] _T_1097; // @[Mux.scala 19:72:@3419.4]
  wire [39:0] _T_1099; // @[Mux.scala 19:72:@3420.4]
  wire [39:0] _T_1101; // @[Mux.scala 19:72:@3421.4]
  wire [39:0] _T_1103; // @[Mux.scala 19:72:@3422.4]
  wire [39:0] _T_1105; // @[Mux.scala 19:72:@3423.4]
  wire [39:0] _T_1107; // @[Mux.scala 19:72:@3424.4]
  wire [39:0] _T_1109; // @[Mux.scala 19:72:@3425.4]
  wire [39:0] _T_1111; // @[Mux.scala 19:72:@3426.4]
  wire [39:0] _T_1113; // @[Mux.scala 19:72:@3427.4]
  wire [39:0] _T_1115; // @[Mux.scala 19:72:@3428.4]
  wire [39:0] _T_1117; // @[Mux.scala 19:72:@3429.4]
  wire [39:0] _T_1119; // @[Mux.scala 19:72:@3430.4]
  wire [39:0] _T_1121; // @[Mux.scala 19:72:@3431.4]
  wire [39:0] _T_1123; // @[Mux.scala 19:72:@3432.4]
  wire [39:0] _T_1125; // @[Mux.scala 19:72:@3433.4]
  wire [63:0] _T_1130; // @[Mux.scala 19:72:@3436.4]
  wire [63:0] _GEN_149; // @[Mux.scala 19:72:@3437.4]
  wire [63:0] _T_1131; // @[Mux.scala 19:72:@3437.4]
  wire [63:0] _GEN_150; // @[Mux.scala 19:72:@3440.4]
  wire [63:0] _T_1134; // @[Mux.scala 19:72:@3440.4]
  wire [63:0] _GEN_151; // @[Mux.scala 19:72:@3441.4]
  wire [63:0] _T_1135; // @[Mux.scala 19:72:@3441.4]
  wire [63:0] _GEN_152; // @[Mux.scala 19:72:@3442.4]
  wire [63:0] _T_1136; // @[Mux.scala 19:72:@3442.4]
  wire [63:0] _GEN_153; // @[Mux.scala 19:72:@3443.4]
  wire [63:0] _T_1137; // @[Mux.scala 19:72:@3443.4]
  wire [63:0] _GEN_154; // @[Mux.scala 19:72:@3444.4]
  wire [63:0] _T_1138; // @[Mux.scala 19:72:@3444.4]
  wire [63:0] _GEN_155; // @[Mux.scala 19:72:@3445.4]
  wire [63:0] _T_1139; // @[Mux.scala 19:72:@3445.4]
  wire [63:0] _GEN_156; // @[Mux.scala 19:72:@3446.4]
  wire [63:0] _T_1140; // @[Mux.scala 19:72:@3446.4]
  wire [63:0] _GEN_157; // @[Mux.scala 19:72:@3447.4]
  wire [63:0] _T_1141; // @[Mux.scala 19:72:@3447.4]
  wire [63:0] _GEN_158; // @[Mux.scala 19:72:@3448.4]
  wire [63:0] _T_1142; // @[Mux.scala 19:72:@3448.4]
  wire [63:0] _GEN_159; // @[Mux.scala 19:72:@3450.4]
  wire [63:0] _T_1144; // @[Mux.scala 19:72:@3450.4]
  wire [63:0] _GEN_160; // @[Mux.scala 19:72:@3451.4]
  wire [63:0] _T_1145; // @[Mux.scala 19:72:@3451.4]
  wire [63:0] _GEN_161; // @[Mux.scala 19:72:@3452.4]
  wire [63:0] _T_1146; // @[Mux.scala 19:72:@3452.4]
  wire [63:0] _GEN_162; // @[Mux.scala 19:72:@3453.4]
  wire [63:0] _T_1147; // @[Mux.scala 19:72:@3453.4]
  wire [63:0] _GEN_163; // @[Mux.scala 19:72:@3454.4]
  wire [63:0] _T_1148; // @[Mux.scala 19:72:@3454.4]
  wire [63:0] _GEN_164; // @[Mux.scala 19:72:@3455.4]
  wire [63:0] _T_1149; // @[Mux.scala 19:72:@3455.4]
  wire [63:0] _GEN_165; // @[Mux.scala 19:72:@3456.4]
  wire [63:0] _T_1150; // @[Mux.scala 19:72:@3456.4]
  wire [63:0] _GEN_166; // @[Mux.scala 19:72:@3457.4]
  wire [63:0] _T_1151; // @[Mux.scala 19:72:@3457.4]
  wire [63:0] _GEN_167; // @[Mux.scala 19:72:@3458.4]
  wire [63:0] _T_1152; // @[Mux.scala 19:72:@3458.4]
  wire [63:0] _GEN_168; // @[Mux.scala 19:72:@3459.4]
  wire [63:0] _T_1153; // @[Mux.scala 19:72:@3459.4]
  wire [63:0] _GEN_169; // @[Mux.scala 19:72:@3460.4]
  wire [63:0] _T_1154; // @[Mux.scala 19:72:@3460.4]
  wire [63:0] _GEN_170; // @[Mux.scala 19:72:@3461.4]
  wire [63:0] _T_1155; // @[Mux.scala 19:72:@3461.4]
  wire [63:0] _GEN_171; // @[Mux.scala 19:72:@3462.4]
  wire [63:0] _T_1156; // @[Mux.scala 19:72:@3462.4]
  wire [63:0] _GEN_172; // @[Mux.scala 19:72:@3463.4]
  wire [63:0] _T_1157; // @[Mux.scala 19:72:@3463.4]
  wire [63:0] _GEN_173; // @[Mux.scala 19:72:@3464.4]
  wire [63:0] _T_1158; // @[Mux.scala 19:72:@3464.4]
  wire [63:0] _GEN_174; // @[Mux.scala 19:72:@3465.4]
  wire [63:0] _T_1159; // @[Mux.scala 19:72:@3465.4]
  wire [63:0] _GEN_175; // @[Mux.scala 19:72:@3466.4]
  wire [63:0] _T_1160; // @[Mux.scala 19:72:@3466.4]
  wire [63:0] _GEN_176; // @[Mux.scala 19:72:@3467.4]
  wire [63:0] _T_1161; // @[Mux.scala 19:72:@3467.4]
  wire [63:0] _GEN_177; // @[Mux.scala 19:72:@3468.4]
  wire [63:0] _T_1162; // @[Mux.scala 19:72:@3468.4]
  wire [63:0] _GEN_178; // @[Mux.scala 19:72:@3469.4]
  wire [63:0] _T_1163; // @[Mux.scala 19:72:@3469.4]
  wire [63:0] _GEN_179; // @[Mux.scala 19:72:@3470.4]
  wire [63:0] _T_1164; // @[Mux.scala 19:72:@3470.4]
  wire [63:0] _GEN_180; // @[Mux.scala 19:72:@3471.4]
  wire [63:0] _T_1165; // @[Mux.scala 19:72:@3471.4]
  wire [63:0] _GEN_181; // @[Mux.scala 19:72:@3472.4]
  wire [63:0] _T_1166; // @[Mux.scala 19:72:@3472.4]
  wire [63:0] _GEN_182; // @[Mux.scala 19:72:@3473.4]
  wire [63:0] _T_1167; // @[Mux.scala 19:72:@3473.4]
  wire [63:0] _GEN_183; // @[Mux.scala 19:72:@3474.4]
  wire [63:0] _T_1168; // @[Mux.scala 19:72:@3474.4]
  wire [63:0] _GEN_184; // @[Mux.scala 19:72:@3475.4]
  wire [63:0] _T_1169; // @[Mux.scala 19:72:@3475.4]
  wire [63:0] _GEN_185; // @[Mux.scala 19:72:@3476.4]
  wire [63:0] _T_1170; // @[Mux.scala 19:72:@3476.4]
  wire [63:0] _GEN_186; // @[Mux.scala 19:72:@3477.4]
  wire [63:0] _T_1171; // @[Mux.scala 19:72:@3477.4]
  wire [63:0] _GEN_187; // @[Mux.scala 19:72:@3478.4]
  wire [63:0] _T_1172; // @[Mux.scala 19:72:@3478.4]
  wire [63:0] _GEN_188; // @[Mux.scala 19:72:@3479.4]
  wire [63:0] _T_1173; // @[Mux.scala 19:72:@3479.4]
  wire [63:0] _GEN_189; // @[Mux.scala 19:72:@3480.4]
  wire [63:0] _T_1174; // @[Mux.scala 19:72:@3480.4]
  wire [63:0] _GEN_190; // @[Mux.scala 19:72:@3481.4]
  wire [63:0] _T_1175; // @[Mux.scala 19:72:@3481.4]
  wire [63:0] _GEN_191; // @[Mux.scala 19:72:@3482.4]
  wire [63:0] _T_1176; // @[Mux.scala 19:72:@3482.4]
  wire [63:0] _GEN_192; // @[Mux.scala 19:72:@3483.4]
  wire [63:0] _T_1177; // @[Mux.scala 19:72:@3483.4]
  wire [63:0] _GEN_193; // @[Mux.scala 19:72:@3484.4]
  wire [63:0] _T_1178; // @[Mux.scala 19:72:@3484.4]
  wire [63:0] _GEN_194; // @[Mux.scala 19:72:@3485.4]
  wire [63:0] _T_1179; // @[Mux.scala 19:72:@3485.4]
  wire [63:0] _GEN_195; // @[Mux.scala 19:72:@3486.4]
  wire [63:0] _T_1180; // @[Mux.scala 19:72:@3486.4]
  wire [63:0] _GEN_196; // @[Mux.scala 19:72:@3487.4]
  wire [63:0] _T_1181; // @[Mux.scala 19:72:@3487.4]
  wire [63:0] _GEN_197; // @[Mux.scala 19:72:@3488.4]
  wire [63:0] _T_1182; // @[Mux.scala 19:72:@3488.4]
  wire [63:0] _GEN_198; // @[Mux.scala 19:72:@3489.4]
  wire [63:0] _T_1183; // @[Mux.scala 19:72:@3489.4]
  wire [63:0] _GEN_199; // @[Mux.scala 19:72:@3490.4]
  wire [63:0] _T_1184; // @[Mux.scala 19:72:@3490.4]
  wire [63:0] _GEN_200; // @[Mux.scala 19:72:@3491.4]
  wire [63:0] _T_1185; // @[Mux.scala 19:72:@3491.4]
  wire [63:0] _GEN_201; // @[Mux.scala 19:72:@3492.4]
  wire [63:0] _T_1186; // @[Mux.scala 19:72:@3492.4]
  wire [63:0] _GEN_202; // @[Mux.scala 19:72:@3493.4]
  wire [63:0] _T_1187; // @[Mux.scala 19:72:@3493.4]
  wire [63:0] _GEN_203; // @[Mux.scala 19:72:@3494.4]
  wire [63:0] _T_1188; // @[Mux.scala 19:72:@3494.4]
  wire [63:0] _GEN_204; // @[Mux.scala 19:72:@3495.4]
  wire [63:0] _T_1189; // @[Mux.scala 19:72:@3495.4]
  wire [63:0] _GEN_205; // @[Mux.scala 19:72:@3496.4]
  wire [63:0] _T_1190; // @[Mux.scala 19:72:@3496.4]
  wire [63:0] _GEN_206; // @[Mux.scala 19:72:@3497.4]
  wire [63:0] _T_1191; // @[Mux.scala 19:72:@3497.4]
  wire [63:0] _GEN_207; // @[Mux.scala 19:72:@3498.4]
  wire [63:0] _T_1192; // @[Mux.scala 19:72:@3498.4]
  wire [63:0] _GEN_208; // @[Mux.scala 19:72:@3499.4]
  wire [63:0] _T_1193; // @[Mux.scala 19:72:@3499.4]
  wire [63:0] _GEN_209; // @[Mux.scala 19:72:@3500.4]
  wire [63:0] _T_1194; // @[Mux.scala 19:72:@3500.4]
  wire [63:0] _GEN_210; // @[Mux.scala 19:72:@3501.4]
  wire [63:0] _T_1195; // @[Mux.scala 19:72:@3501.4]
  wire [63:0] _GEN_211; // @[Mux.scala 19:72:@3502.4]
  wire [63:0] _T_1196; // @[Mux.scala 19:72:@3502.4]
  wire [63:0] _GEN_212; // @[Mux.scala 19:72:@3503.4]
  wire [63:0] _T_1197; // @[Mux.scala 19:72:@3503.4]
  wire [63:0] _GEN_213; // @[Mux.scala 19:72:@3504.4]
  wire [63:0] _T_1198; // @[Mux.scala 19:72:@3504.4]
  wire [63:0] _GEN_214; // @[Mux.scala 19:72:@3505.4]
  wire [63:0] _T_1199; // @[Mux.scala 19:72:@3505.4]
  wire [63:0] _GEN_215; // @[Mux.scala 19:72:@3506.4]
  wire [63:0] _T_1200; // @[Mux.scala 19:72:@3506.4]
  wire [63:0] _GEN_216; // @[Mux.scala 19:72:@3507.4]
  wire [63:0] _T_1201; // @[Mux.scala 19:72:@3507.4]
  wire [63:0] _GEN_217; // @[Mux.scala 19:72:@3508.4]
  wire [63:0] _T_1202; // @[Mux.scala 19:72:@3508.4]
  wire [63:0] _GEN_218; // @[Mux.scala 19:72:@3509.4]
  wire [63:0] _T_1203; // @[Mux.scala 19:72:@3509.4]
  wire [63:0] _GEN_219; // @[Mux.scala 19:72:@3510.4]
  wire [63:0] _T_1204; // @[Mux.scala 19:72:@3510.4]
  wire [63:0] _GEN_220; // @[Mux.scala 19:72:@3511.4]
  wire [63:0] _T_1205; // @[Mux.scala 19:72:@3511.4]
  wire [63:0] _GEN_221; // @[Mux.scala 19:72:@3512.4]
  wire [63:0] _T_1206; // @[Mux.scala 19:72:@3512.4]
  wire [63:0] _GEN_222; // @[Mux.scala 19:72:@3513.4]
  wire [63:0] _T_1207; // @[Mux.scala 19:72:@3513.4]
  wire [63:0] _GEN_223; // @[Mux.scala 19:72:@3514.4]
  wire [63:0] _T_1208; // @[Mux.scala 19:72:@3514.4]
  wire [63:0] _GEN_224; // @[Mux.scala 19:72:@3515.4]
  wire [63:0] _T_1209; // @[Mux.scala 19:72:@3515.4]
  wire  _T_1220; // @[CSR.scala 245:39:@3528.8]
  wire  _T_1222; // @[CSR.scala 245:39:@3532.8]
  wire  _GEN_17; // @[CSR.scala 244:39:@3522.6]
  wire  _GEN_18; // @[CSR.scala 244:39:@3522.6]
  wire [15:0] _T_1233; // @[:@3551.8 :@3552.8]
  wire  _T_1235; // @[CSR.scala 250:35:@3555.8]
  wire  _T_1237; // @[CSR.scala 250:35:@3559.8]
  wire  _GEN_19; // @[CSR.scala 249:35:@3549.6]
  wire  _GEN_20; // @[CSR.scala 253:35:@3569.6]
  wire  _GEN_21; // @[CSR.scala 253:35:@3569.6]
  wire [7:0] _T_1253; // @[CSR.scala 277:47:@3591.8]
  wire [31:0] _T_1254; // @[CSR.scala 277:72:@3592.8]
  wire [39:0] _T_1255; // @[Cat.scala 30:58:@3593.8]
  wire [40:0] _GEN_22; // @[CSR.scala 277:29:@3590.6]
  wire [7:0] _T_1256; // @[CSR.scala 278:45:@3597.8]
  wire [39:0] _T_1257; // @[Cat.scala 30:58:@3598.8]
  wire [40:0] _GEN_23; // @[CSR.scala 278:29:@3596.6]
  wire [31:0] _T_1259; // @[CSR.scala 277:72:@3603.8]
  wire [39:0] _T_1260; // @[Cat.scala 30:58:@3604.8]
  wire [40:0] _GEN_24; // @[CSR.scala 277:29:@3601.6]
  wire [7:0] _T_1261; // @[CSR.scala 278:45:@3608.8]
  wire [39:0] _T_1262; // @[Cat.scala 30:58:@3609.8]
  wire [40:0] _GEN_25; // @[CSR.scala 278:29:@3607.6]
  wire [31:0] _T_1264; // @[CSR.scala 277:72:@3614.8]
  wire [39:0] _T_1265; // @[Cat.scala 30:58:@3615.8]
  wire [40:0] _GEN_26; // @[CSR.scala 277:29:@3612.6]
  wire [7:0] _T_1266; // @[CSR.scala 278:45:@3619.8]
  wire [39:0] _T_1267; // @[Cat.scala 30:58:@3620.8]
  wire [40:0] _GEN_27; // @[CSR.scala 278:29:@3618.6]
  wire [31:0] _T_1269; // @[CSR.scala 277:72:@3625.8]
  wire [39:0] _T_1270; // @[Cat.scala 30:58:@3626.8]
  wire [40:0] _GEN_28; // @[CSR.scala 277:29:@3623.6]
  wire [7:0] _T_1271; // @[CSR.scala 278:45:@3630.8]
  wire [39:0] _T_1272; // @[Cat.scala 30:58:@3631.8]
  wire [40:0] _GEN_29; // @[CSR.scala 278:29:@3629.6]
  wire [31:0] _T_1274; // @[CSR.scala 277:72:@3636.8]
  wire [39:0] _T_1275; // @[Cat.scala 30:58:@3637.8]
  wire [40:0] _GEN_30; // @[CSR.scala 277:29:@3634.6]
  wire [7:0] _T_1276; // @[CSR.scala 278:45:@3641.8]
  wire [39:0] _T_1277; // @[Cat.scala 30:58:@3642.8]
  wire [40:0] _GEN_31; // @[CSR.scala 278:29:@3640.6]
  wire [31:0] _T_1279; // @[CSR.scala 277:72:@3647.8]
  wire [39:0] _T_1280; // @[Cat.scala 30:58:@3648.8]
  wire [40:0] _GEN_32; // @[CSR.scala 277:29:@3645.6]
  wire [7:0] _T_1281; // @[CSR.scala 278:45:@3652.8]
  wire [39:0] _T_1282; // @[Cat.scala 30:58:@3653.8]
  wire [40:0] _GEN_33; // @[CSR.scala 278:29:@3651.6]
  wire [31:0] _T_1284; // @[CSR.scala 277:72:@3658.8]
  wire [39:0] _T_1285; // @[Cat.scala 30:58:@3659.8]
  wire [40:0] _GEN_34; // @[CSR.scala 277:29:@3656.6]
  wire [7:0] _T_1286; // @[CSR.scala 278:45:@3663.8]
  wire [39:0] _T_1287; // @[Cat.scala 30:58:@3664.8]
  wire [40:0] _GEN_35; // @[CSR.scala 278:29:@3662.6]
  wire [31:0] _T_1289; // @[CSR.scala 277:72:@3669.8]
  wire [39:0] _T_1290; // @[Cat.scala 30:58:@3670.8]
  wire [40:0] _GEN_36; // @[CSR.scala 277:29:@3667.6]
  wire [7:0] _T_1291; // @[CSR.scala 278:45:@3674.8]
  wire [39:0] _T_1292; // @[Cat.scala 30:58:@3675.8]
  wire [40:0] _GEN_37; // @[CSR.scala 278:29:@3673.6]
  wire [31:0] _T_1294; // @[CSR.scala 277:72:@3680.8]
  wire [39:0] _T_1295; // @[Cat.scala 30:58:@3681.8]
  wire [40:0] _GEN_38; // @[CSR.scala 277:29:@3678.6]
  wire [7:0] _T_1296; // @[CSR.scala 278:45:@3685.8]
  wire [39:0] _T_1297; // @[Cat.scala 30:58:@3686.8]
  wire [40:0] _GEN_39; // @[CSR.scala 278:29:@3684.6]
  wire [31:0] _T_1299; // @[CSR.scala 277:72:@3691.8]
  wire [39:0] _T_1300; // @[Cat.scala 30:58:@3692.8]
  wire [40:0] _GEN_40; // @[CSR.scala 277:29:@3689.6]
  wire [7:0] _T_1301; // @[CSR.scala 278:45:@3696.8]
  wire [39:0] _T_1302; // @[Cat.scala 30:58:@3697.8]
  wire [40:0] _GEN_41; // @[CSR.scala 278:29:@3695.6]
  wire [31:0] _T_1304; // @[CSR.scala 277:72:@3702.8]
  wire [39:0] _T_1305; // @[Cat.scala 30:58:@3703.8]
  wire [40:0] _GEN_42; // @[CSR.scala 277:29:@3700.6]
  wire [7:0] _T_1306; // @[CSR.scala 278:45:@3707.8]
  wire [39:0] _T_1307; // @[Cat.scala 30:58:@3708.8]
  wire [40:0] _GEN_43; // @[CSR.scala 278:29:@3706.6]
  wire [31:0] _T_1309; // @[CSR.scala 277:72:@3713.8]
  wire [39:0] _T_1310; // @[Cat.scala 30:58:@3714.8]
  wire [40:0] _GEN_44; // @[CSR.scala 277:29:@3711.6]
  wire [7:0] _T_1311; // @[CSR.scala 278:45:@3718.8]
  wire [39:0] _T_1312; // @[Cat.scala 30:58:@3719.8]
  wire [40:0] _GEN_45; // @[CSR.scala 278:29:@3717.6]
  wire [31:0] _T_1314; // @[CSR.scala 277:72:@3724.8]
  wire [39:0] _T_1315; // @[Cat.scala 30:58:@3725.8]
  wire [40:0] _GEN_46; // @[CSR.scala 277:29:@3722.6]
  wire [7:0] _T_1316; // @[CSR.scala 278:45:@3729.8]
  wire [39:0] _T_1317; // @[Cat.scala 30:58:@3730.8]
  wire [40:0] _GEN_47; // @[CSR.scala 278:29:@3728.6]
  wire [31:0] _T_1319; // @[CSR.scala 277:72:@3735.8]
  wire [39:0] _T_1320; // @[Cat.scala 30:58:@3736.8]
  wire [40:0] _GEN_48; // @[CSR.scala 277:29:@3733.6]
  wire [7:0] _T_1321; // @[CSR.scala 278:45:@3740.8]
  wire [39:0] _T_1322; // @[Cat.scala 30:58:@3741.8]
  wire [40:0] _GEN_49; // @[CSR.scala 278:29:@3739.6]
  wire [31:0] _T_1324; // @[CSR.scala 277:72:@3746.8]
  wire [39:0] _T_1325; // @[Cat.scala 30:58:@3747.8]
  wire [40:0] _GEN_50; // @[CSR.scala 277:29:@3744.6]
  wire [7:0] _T_1326; // @[CSR.scala 278:45:@3751.8]
  wire [39:0] _T_1327; // @[Cat.scala 30:58:@3752.8]
  wire [40:0] _GEN_51; // @[CSR.scala 278:29:@3750.6]
  wire [31:0] _T_1329; // @[CSR.scala 277:72:@3757.8]
  wire [39:0] _T_1330; // @[Cat.scala 30:58:@3758.8]
  wire [40:0] _GEN_52; // @[CSR.scala 277:29:@3755.6]
  wire [7:0] _T_1331; // @[CSR.scala 278:45:@3762.8]
  wire [39:0] _T_1332; // @[Cat.scala 30:58:@3763.8]
  wire [40:0] _GEN_53; // @[CSR.scala 278:29:@3761.6]
  wire [31:0] _T_1334; // @[CSR.scala 277:72:@3768.8]
  wire [39:0] _T_1335; // @[Cat.scala 30:58:@3769.8]
  wire [40:0] _GEN_54; // @[CSR.scala 277:29:@3766.6]
  wire [7:0] _T_1336; // @[CSR.scala 278:45:@3773.8]
  wire [39:0] _T_1337; // @[Cat.scala 30:58:@3774.8]
  wire [40:0] _GEN_55; // @[CSR.scala 278:29:@3772.6]
  wire [31:0] _T_1339; // @[CSR.scala 277:72:@3779.8]
  wire [39:0] _T_1340; // @[Cat.scala 30:58:@3780.8]
  wire [40:0] _GEN_56; // @[CSR.scala 277:29:@3777.6]
  wire [7:0] _T_1341; // @[CSR.scala 278:45:@3784.8]
  wire [39:0] _T_1342; // @[Cat.scala 30:58:@3785.8]
  wire [40:0] _GEN_57; // @[CSR.scala 278:29:@3783.6]
  wire [31:0] _T_1344; // @[CSR.scala 277:72:@3790.8]
  wire [39:0] _T_1345; // @[Cat.scala 30:58:@3791.8]
  wire [40:0] _GEN_58; // @[CSR.scala 277:29:@3788.6]
  wire [7:0] _T_1346; // @[CSR.scala 278:45:@3795.8]
  wire [39:0] _T_1347; // @[Cat.scala 30:58:@3796.8]
  wire [40:0] _GEN_59; // @[CSR.scala 278:29:@3794.6]
  wire [31:0] _T_1349; // @[CSR.scala 277:72:@3801.8]
  wire [39:0] _T_1350; // @[Cat.scala 30:58:@3802.8]
  wire [40:0] _GEN_60; // @[CSR.scala 277:29:@3799.6]
  wire [7:0] _T_1351; // @[CSR.scala 278:45:@3806.8]
  wire [39:0] _T_1352; // @[Cat.scala 30:58:@3807.8]
  wire [40:0] _GEN_61; // @[CSR.scala 278:29:@3805.6]
  wire [31:0] _T_1354; // @[CSR.scala 277:72:@3812.8]
  wire [39:0] _T_1355; // @[Cat.scala 30:58:@3813.8]
  wire [40:0] _GEN_62; // @[CSR.scala 277:29:@3810.6]
  wire [7:0] _T_1356; // @[CSR.scala 278:45:@3817.8]
  wire [39:0] _T_1357; // @[Cat.scala 30:58:@3818.8]
  wire [40:0] _GEN_63; // @[CSR.scala 278:29:@3816.6]
  wire [31:0] _T_1359; // @[CSR.scala 277:72:@3823.8]
  wire [39:0] _T_1360; // @[Cat.scala 30:58:@3824.8]
  wire [40:0] _GEN_64; // @[CSR.scala 277:29:@3821.6]
  wire [7:0] _T_1361; // @[CSR.scala 278:45:@3828.8]
  wire [39:0] _T_1362; // @[Cat.scala 30:58:@3829.8]
  wire [40:0] _GEN_65; // @[CSR.scala 278:29:@3827.6]
  wire [31:0] _T_1364; // @[CSR.scala 277:72:@3834.8]
  wire [39:0] _T_1365; // @[Cat.scala 30:58:@3835.8]
  wire [40:0] _GEN_66; // @[CSR.scala 277:29:@3832.6]
  wire [7:0] _T_1366; // @[CSR.scala 278:45:@3839.8]
  wire [39:0] _T_1367; // @[Cat.scala 30:58:@3840.8]
  wire [40:0] _GEN_67; // @[CSR.scala 278:29:@3838.6]
  wire [31:0] _T_1369; // @[CSR.scala 277:72:@3845.8]
  wire [39:0] _T_1370; // @[Cat.scala 30:58:@3846.8]
  wire [40:0] _GEN_68; // @[CSR.scala 277:29:@3843.6]
  wire [7:0] _T_1371; // @[CSR.scala 278:45:@3850.8]
  wire [39:0] _T_1372; // @[Cat.scala 30:58:@3851.8]
  wire [40:0] _GEN_69; // @[CSR.scala 278:29:@3849.6]
  wire [31:0] _T_1374; // @[CSR.scala 277:72:@3856.8]
  wire [39:0] _T_1375; // @[Cat.scala 30:58:@3857.8]
  wire [40:0] _GEN_70; // @[CSR.scala 277:29:@3854.6]
  wire [7:0] _T_1376; // @[CSR.scala 278:45:@3861.8]
  wire [39:0] _T_1377; // @[Cat.scala 30:58:@3862.8]
  wire [40:0] _GEN_71; // @[CSR.scala 278:29:@3860.6]
  wire [31:0] _T_1379; // @[CSR.scala 277:72:@3867.8]
  wire [39:0] _T_1380; // @[Cat.scala 30:58:@3868.8]
  wire [40:0] _GEN_72; // @[CSR.scala 277:29:@3865.6]
  wire [7:0] _T_1381; // @[CSR.scala 278:45:@3872.8]
  wire [39:0] _T_1382; // @[Cat.scala 30:58:@3873.8]
  wire [40:0] _GEN_73; // @[CSR.scala 278:29:@3871.6]
  wire [31:0] _T_1384; // @[CSR.scala 277:72:@3878.8]
  wire [39:0] _T_1385; // @[Cat.scala 30:58:@3879.8]
  wire [40:0] _GEN_74; // @[CSR.scala 277:29:@3876.6]
  wire [7:0] _T_1386; // @[CSR.scala 278:45:@3883.8]
  wire [39:0] _T_1387; // @[Cat.scala 30:58:@3884.8]
  wire [40:0] _GEN_75; // @[CSR.scala 278:29:@3882.6]
  wire [31:0] _T_1389; // @[CSR.scala 277:72:@3889.8]
  wire [39:0] _T_1390; // @[Cat.scala 30:58:@3890.8]
  wire [40:0] _GEN_76; // @[CSR.scala 277:29:@3887.6]
  wire [7:0] _T_1391; // @[CSR.scala 278:45:@3894.8]
  wire [39:0] _T_1392; // @[Cat.scala 30:58:@3895.8]
  wire [40:0] _GEN_77; // @[CSR.scala 278:29:@3893.6]
  wire [31:0] _T_1394; // @[CSR.scala 277:72:@3900.8]
  wire [39:0] _T_1395; // @[Cat.scala 30:58:@3901.8]
  wire [40:0] _GEN_78; // @[CSR.scala 277:29:@3898.6]
  wire [7:0] _T_1396; // @[CSR.scala 278:45:@3905.8]
  wire [39:0] _T_1397; // @[Cat.scala 30:58:@3906.8]
  wire [40:0] _GEN_79; // @[CSR.scala 278:29:@3904.6]
  wire [31:0] _T_1399; // @[CSR.scala 277:72:@3911.8]
  wire [39:0] _T_1400; // @[Cat.scala 30:58:@3912.8]
  wire [40:0] _GEN_80; // @[CSR.scala 277:29:@3909.6]
  wire [7:0] _T_1401; // @[CSR.scala 278:45:@3916.8]
  wire [39:0] _T_1402; // @[Cat.scala 30:58:@3917.8]
  wire [40:0] _GEN_81; // @[CSR.scala 278:29:@3915.6]
  wire [31:0] _T_1404; // @[CSR.scala 277:72:@3922.8]
  wire [39:0] _T_1405; // @[Cat.scala 30:58:@3923.8]
  wire [40:0] _GEN_82; // @[CSR.scala 277:29:@3920.6]
  wire [7:0] _T_1406; // @[CSR.scala 278:45:@3927.8]
  wire [39:0] _T_1407; // @[Cat.scala 30:58:@3928.8]
  wire [40:0] _GEN_83; // @[CSR.scala 278:29:@3926.6]
  wire [31:0] _T_1409; // @[CSR.scala 277:72:@3933.8]
  wire [39:0] _T_1410; // @[Cat.scala 30:58:@3934.8]
  wire [40:0] _GEN_84; // @[CSR.scala 277:29:@3931.6]
  wire [7:0] _T_1411; // @[CSR.scala 278:45:@3938.8]
  wire [39:0] _T_1412; // @[Cat.scala 30:58:@3939.8]
  wire [40:0] _GEN_85; // @[CSR.scala 278:29:@3937.6]
  wire [31:0] _T_1414; // @[CSR.scala 277:72:@3944.8]
  wire [63:0] _T_1415; // @[Cat.scala 30:58:@3945.8]
  wire [57:0] _T_1416; // @[Util.scala 133:28:@3947.8]
  wire [63:0] _GEN_86; // @[CSR.scala 277:29:@3942.6]
  wire [57:0] _GEN_87; // @[CSR.scala 277:29:@3942.6]
  wire [31:0] _T_1417; // @[CSR.scala 278:45:@3951.8]
  wire [63:0] _T_1418; // @[Cat.scala 30:58:@3952.8]
  wire [57:0] _T_1419; // @[Util.scala 133:28:@3954.8]
  wire [63:0] _GEN_88; // @[CSR.scala 278:29:@3950.6]
  wire [57:0] _GEN_89; // @[CSR.scala 278:29:@3950.6]
  wire [31:0] _T_1421; // @[CSR.scala 277:72:@3959.8]
  wire [63:0] _T_1422; // @[Cat.scala 30:58:@3960.8]
  wire [57:0] _T_1423; // @[Util.scala 133:28:@3962.8]
  wire [63:0] _GEN_90; // @[CSR.scala 277:29:@3957.6]
  wire [57:0] _GEN_91; // @[CSR.scala 277:29:@3957.6]
  wire [31:0] _T_1424; // @[CSR.scala 278:45:@3966.8]
  wire [63:0] _T_1425; // @[Cat.scala 30:58:@3967.8]
  wire [57:0] _T_1426; // @[Util.scala 133:28:@3969.8]
  wire [63:0] _GEN_92; // @[CSR.scala 278:29:@3965.6]
  wire [57:0] _GEN_93; // @[CSR.scala 278:29:@3965.6]
  wire [31:0] _GEN_94; // @[CSR.scala 265:40:@3972.6]
  wire [31:0] _T_1429; // @[CSR.scala 267:78:@3977.8]
  wire [34:0] _GEN_225; // @[CSR.scala 267:86:@3978.8]
  wire [34:0] _T_1431; // @[CSR.scala 267:86:@3978.8]
  wire [34:0] _GEN_95; // @[CSR.scala 267:40:@3975.6]
  wire [31:0] _GEN_96; // @[CSR.scala 268:40:@3981.6]
  wire [31:0] _T_1433; // @[CSR.scala 269:62:@3985.8]
  wire [31:0] _GEN_97; // @[CSR.scala 269:40:@3984.6]
  wire [31:0] _GEN_98; // @[CSR.scala 270:40:@3988.6]
  wire [31:0] _GEN_99; // @[CSR.scala 271:42:@3992.6]
  wire  _GEN_100; // @[CSR.scala 242:14:@3521.4]
  wire  _GEN_101; // @[CSR.scala 242:14:@3521.4]
  wire  _GEN_102; // @[CSR.scala 242:14:@3521.4]
  wire  _GEN_103; // @[CSR.scala 242:14:@3521.4]
  wire  _GEN_104; // @[CSR.scala 242:14:@3521.4]
  wire [40:0] _GEN_105; // @[CSR.scala 242:14:@3521.4]
  wire [40:0] _GEN_106; // @[CSR.scala 242:14:@3521.4]
  wire [40:0] _GEN_107; // @[CSR.scala 242:14:@3521.4]
  wire [40:0] _GEN_108; // @[CSR.scala 242:14:@3521.4]
  wire [40:0] _GEN_109; // @[CSR.scala 242:14:@3521.4]
  wire [40:0] _GEN_110; // @[CSR.scala 242:14:@3521.4]
  wire [40:0] _GEN_111; // @[CSR.scala 242:14:@3521.4]
  wire [40:0] _GEN_112; // @[CSR.scala 242:14:@3521.4]
  wire [40:0] _GEN_113; // @[CSR.scala 242:14:@3521.4]
  wire [40:0] _GEN_114; // @[CSR.scala 242:14:@3521.4]
  wire [40:0] _GEN_115; // @[CSR.scala 242:14:@3521.4]
  wire [40:0] _GEN_116; // @[CSR.scala 242:14:@3521.4]
  wire [40:0] _GEN_117; // @[CSR.scala 242:14:@3521.4]
  wire [40:0] _GEN_118; // @[CSR.scala 242:14:@3521.4]
  wire [40:0] _GEN_119; // @[CSR.scala 242:14:@3521.4]
  wire [40:0] _GEN_120; // @[CSR.scala 242:14:@3521.4]
  wire [40:0] _GEN_121; // @[CSR.scala 242:14:@3521.4]
  wire [40:0] _GEN_122; // @[CSR.scala 242:14:@3521.4]
  wire [40:0] _GEN_123; // @[CSR.scala 242:14:@3521.4]
  wire [40:0] _GEN_124; // @[CSR.scala 242:14:@3521.4]
  wire [40:0] _GEN_125; // @[CSR.scala 242:14:@3521.4]
  wire [40:0] _GEN_126; // @[CSR.scala 242:14:@3521.4]
  wire [40:0] _GEN_127; // @[CSR.scala 242:14:@3521.4]
  wire [40:0] _GEN_128; // @[CSR.scala 242:14:@3521.4]
  wire [40:0] _GEN_129; // @[CSR.scala 242:14:@3521.4]
  wire [40:0] _GEN_130; // @[CSR.scala 242:14:@3521.4]
  wire [40:0] _GEN_131; // @[CSR.scala 242:14:@3521.4]
  wire [40:0] _GEN_132; // @[CSR.scala 242:14:@3521.4]
  wire [40:0] _GEN_133; // @[CSR.scala 242:14:@3521.4]
  wire [40:0] _GEN_134; // @[CSR.scala 242:14:@3521.4]
  wire [40:0] _GEN_135; // @[CSR.scala 242:14:@3521.4]
  wire [40:0] _GEN_136; // @[CSR.scala 242:14:@3521.4]
  wire [63:0] _GEN_137; // @[CSR.scala 242:14:@3521.4]
  wire [57:0] _GEN_138; // @[CSR.scala 242:14:@3521.4]
  wire [63:0] _GEN_139; // @[CSR.scala 242:14:@3521.4]
  wire [57:0] _GEN_140; // @[CSR.scala 242:14:@3521.4]
  wire [34:0] _GEN_142; // @[CSR.scala 242:14:@3521.4]
  assign _T_241 = _T_240 + 6'h1; // @[Util.scala 113:33:@2767.4]
  assign _T_245 = _T_241[6]; // @[Util.scala 118:20:@2770.4]
  assign _T_247 = _T_244 + 58'h1; // @[Util.scala 118:43:@2772.6]
  assign _T_248 = _T_244 + 58'h1; // @[Util.scala 118:43:@2773.6]
  assign _GEN_0 = _T_245 ? _T_248 : _T_244; // @[Util.scala 118:34:@2771.4]
  assign _T_249 = {_T_244,_T_240}; // @[Cat.scala 30:58:@2776.4]
  assign _GEN_147 = {{4'd0}, io_retire}; // @[Util.scala 113:33:@2778.4]
  assign _T_253 = _T_252 + _GEN_147; // @[Util.scala 113:33:@2778.4]
  assign _T_257 = _T_253[6]; // @[Util.scala 118:20:@2781.4]
  assign _T_259 = _T_256 + 58'h1; // @[Util.scala 118:43:@2783.6]
  assign _T_260 = _T_256 + 58'h1; // @[Util.scala 118:43:@2784.6]
  assign _GEN_1 = _T_257 ? _T_260 : _T_256; // @[Util.scala 118:34:@2782.4]
  assign _T_261 = {_T_256,_T_252}; // @[Cat.scala 30:58:@2787.4]
  assign _T_265 = {{1'd0}, _T_264}; // @[Util.scala 113:33:@2790.4]
  assign _T_268 = {{1'd0}, _T_267}; // @[Util.scala 113:33:@2793.4]
  assign _T_271 = {{1'd0}, _T_270}; // @[Util.scala 113:33:@2796.4]
  assign _T_274 = {{1'd0}, _T_273}; // @[Util.scala 113:33:@2799.4]
  assign _T_277 = {{1'd0}, _T_276}; // @[Util.scala 113:33:@2802.4]
  assign _T_280 = {{1'd0}, _T_279}; // @[Util.scala 113:33:@2805.4]
  assign _T_283 = {{1'd0}, _T_282}; // @[Util.scala 113:33:@2808.4]
  assign _T_286 = {{1'd0}, _T_285}; // @[Util.scala 113:33:@2811.4]
  assign _T_289 = {{1'd0}, _T_288}; // @[Util.scala 113:33:@2814.4]
  assign _T_292 = {{1'd0}, _T_291}; // @[Util.scala 113:33:@2817.4]
  assign _T_295 = {{1'd0}, _T_294}; // @[Util.scala 113:33:@2820.4]
  assign _T_298 = {{1'd0}, _T_297}; // @[Util.scala 113:33:@2823.4]
  assign _T_301 = {{1'd0}, _T_300}; // @[Util.scala 113:33:@2826.4]
  assign _T_304 = {{1'd0}, _T_303}; // @[Util.scala 113:33:@2829.4]
  assign _T_307 = {{1'd0}, _T_306}; // @[Util.scala 113:33:@2832.4]
  assign _T_310 = {{1'd0}, _T_309}; // @[Util.scala 113:33:@2835.4]
  assign _T_313 = {{1'd0}, _T_312}; // @[Util.scala 113:33:@2838.4]
  assign _T_316 = {{1'd0}, _T_315}; // @[Util.scala 113:33:@2841.4]
  assign _T_319 = {{1'd0}, _T_318}; // @[Util.scala 113:33:@2844.4]
  assign _T_322 = {{1'd0}, _T_321}; // @[Util.scala 113:33:@2847.4]
  assign _T_325 = {{1'd0}, _T_324}; // @[Util.scala 113:33:@2850.4]
  assign _T_328 = {{1'd0}, _T_327}; // @[Util.scala 113:33:@2853.4]
  assign _T_331 = {{1'd0}, _T_330}; // @[Util.scala 113:33:@2856.4]
  assign _T_334 = {{1'd0}, _T_333}; // @[Util.scala 113:33:@2859.4]
  assign _T_337 = {{1'd0}, _T_336}; // @[Util.scala 113:33:@2862.4]
  assign _T_340 = {{1'd0}, _T_339}; // @[Util.scala 113:33:@2865.4]
  assign _T_343 = {{1'd0}, _T_342}; // @[Util.scala 113:33:@2868.4]
  assign _T_346 = {{1'd0}, _T_345}; // @[Util.scala 113:33:@2871.4]
  assign _T_349 = {{1'd0}, _T_348}; // @[Util.scala 113:33:@2874.4]
  assign _T_352 = {{1'd0}, _T_351}; // @[Util.scala 113:33:@2877.4]
  assign _T_355 = {{1'd0}, _T_354}; // @[Util.scala 113:33:@2880.4]
  assign _T_358 = {{1'd0}, _T_357}; // @[Util.scala 113:33:@2883.4]
  assign system_insn = io_rw_cmd == 3'h4; // @[CSR.scala 137:31:@2974.4]
  assign _T_446 = io_rw_cmd != 3'h0; // @[CSR.scala 138:27:@2975.4]
  assign _T_448 = system_insn == 1'h0; // @[CSR.scala 138:40:@2976.4]
  assign cpu_ren = _T_446 & _T_448; // @[CSR.scala 138:37:@2977.4]
  assign read_mstatus = {io_status_prv,io_status_unimp5,io_status_mprv,io_status_unimp4,io_status_mpp,io_status_unimp3,io_status_mpie,io_status_unimp2,io_status_mie,io_status_unimp1}; // @[CSR.scala 140:32:@2986.4]
  assign _T_468 = {5'h0,3'h0,reg_mip_mtip,3'h0,reg_mip_msip,3'h0}; // @[CSR.scala 156:25:@2992.4]
  assign _T_474 = {5'h0,3'h0,reg_mie_mtip,3'h0,reg_mie_msip,3'h0}; // @[CSR.scala 157:25:@2998.4]
  assign _T_478 = io_rw_addr == 12'hb00; // @[CSR.scala 177:73:@2999.4]
  assign _T_480 = io_rw_addr == 12'hb02; // @[CSR.scala 177:73:@3000.4]
  assign _T_482 = io_rw_addr == 12'hf13; // @[CSR.scala 177:73:@3001.4]
  assign _T_488 = io_rw_addr == 12'h301; // @[CSR.scala 177:73:@3004.4]
  assign _T_490 = io_rw_addr == 12'h300; // @[CSR.scala 177:73:@3005.4]
  assign _T_492 = io_rw_addr == 12'h305; // @[CSR.scala 177:73:@3006.4]
  assign _T_494 = io_rw_addr == 12'h344; // @[CSR.scala 177:73:@3007.4]
  assign _T_496 = io_rw_addr == 12'h304; // @[CSR.scala 177:73:@3008.4]
  assign _T_498 = io_rw_addr == 12'h340; // @[CSR.scala 177:73:@3009.4]
  assign _T_500 = io_rw_addr == 12'h341; // @[CSR.scala 177:73:@3010.4]
  assign _T_502 = io_rw_addr == 12'h343; // @[CSR.scala 177:73:@3011.4]
  assign _T_504 = io_rw_addr == 12'h342; // @[CSR.scala 177:73:@3012.4]
  assign _T_508 = io_rw_addr == 12'h7b2; // @[CSR.scala 177:73:@3014.4]
  assign _T_510 = io_rw_addr == 12'h302; // @[CSR.scala 177:73:@3015.4]
  assign _T_512 = io_rw_addr == 12'hb03; // @[CSR.scala 177:73:@3016.4]
  assign _T_514 = io_rw_addr == 12'hb83; // @[CSR.scala 177:73:@3017.4]
  assign _T_516 = io_rw_addr == 12'hb04; // @[CSR.scala 177:73:@3018.4]
  assign _T_518 = io_rw_addr == 12'hb84; // @[CSR.scala 177:73:@3019.4]
  assign _T_520 = io_rw_addr == 12'hb05; // @[CSR.scala 177:73:@3020.4]
  assign _T_522 = io_rw_addr == 12'hb85; // @[CSR.scala 177:73:@3021.4]
  assign _T_524 = io_rw_addr == 12'hb06; // @[CSR.scala 177:73:@3022.4]
  assign _T_526 = io_rw_addr == 12'hb86; // @[CSR.scala 177:73:@3023.4]
  assign _T_528 = io_rw_addr == 12'hb07; // @[CSR.scala 177:73:@3024.4]
  assign _T_530 = io_rw_addr == 12'hb87; // @[CSR.scala 177:73:@3025.4]
  assign _T_532 = io_rw_addr == 12'hb08; // @[CSR.scala 177:73:@3026.4]
  assign _T_534 = io_rw_addr == 12'hb88; // @[CSR.scala 177:73:@3027.4]
  assign _T_536 = io_rw_addr == 12'hb09; // @[CSR.scala 177:73:@3028.4]
  assign _T_538 = io_rw_addr == 12'hb89; // @[CSR.scala 177:73:@3029.4]
  assign _T_540 = io_rw_addr == 12'hb0a; // @[CSR.scala 177:73:@3030.4]
  assign _T_542 = io_rw_addr == 12'hb8a; // @[CSR.scala 177:73:@3031.4]
  assign _T_544 = io_rw_addr == 12'hb0b; // @[CSR.scala 177:73:@3032.4]
  assign _T_546 = io_rw_addr == 12'hb8b; // @[CSR.scala 177:73:@3033.4]
  assign _T_548 = io_rw_addr == 12'hb0c; // @[CSR.scala 177:73:@3034.4]
  assign _T_550 = io_rw_addr == 12'hb8c; // @[CSR.scala 177:73:@3035.4]
  assign _T_552 = io_rw_addr == 12'hb0d; // @[CSR.scala 177:73:@3036.4]
  assign _T_554 = io_rw_addr == 12'hb8d; // @[CSR.scala 177:73:@3037.4]
  assign _T_556 = io_rw_addr == 12'hb0e; // @[CSR.scala 177:73:@3038.4]
  assign _T_558 = io_rw_addr == 12'hb8e; // @[CSR.scala 177:73:@3039.4]
  assign _T_560 = io_rw_addr == 12'hb0f; // @[CSR.scala 177:73:@3040.4]
  assign _T_562 = io_rw_addr == 12'hb8f; // @[CSR.scala 177:73:@3041.4]
  assign _T_564 = io_rw_addr == 12'hb10; // @[CSR.scala 177:73:@3042.4]
  assign _T_566 = io_rw_addr == 12'hb90; // @[CSR.scala 177:73:@3043.4]
  assign _T_568 = io_rw_addr == 12'hb11; // @[CSR.scala 177:73:@3044.4]
  assign _T_570 = io_rw_addr == 12'hb91; // @[CSR.scala 177:73:@3045.4]
  assign _T_572 = io_rw_addr == 12'hb12; // @[CSR.scala 177:73:@3046.4]
  assign _T_574 = io_rw_addr == 12'hb92; // @[CSR.scala 177:73:@3047.4]
  assign _T_576 = io_rw_addr == 12'hb13; // @[CSR.scala 177:73:@3048.4]
  assign _T_578 = io_rw_addr == 12'hb93; // @[CSR.scala 177:73:@3049.4]
  assign _T_580 = io_rw_addr == 12'hb14; // @[CSR.scala 177:73:@3050.4]
  assign _T_582 = io_rw_addr == 12'hb94; // @[CSR.scala 177:73:@3051.4]
  assign _T_584 = io_rw_addr == 12'hb15; // @[CSR.scala 177:73:@3052.4]
  assign _T_586 = io_rw_addr == 12'hb95; // @[CSR.scala 177:73:@3053.4]
  assign _T_588 = io_rw_addr == 12'hb16; // @[CSR.scala 177:73:@3054.4]
  assign _T_590 = io_rw_addr == 12'hb96; // @[CSR.scala 177:73:@3055.4]
  assign _T_592 = io_rw_addr == 12'hb17; // @[CSR.scala 177:73:@3056.4]
  assign _T_594 = io_rw_addr == 12'hb97; // @[CSR.scala 177:73:@3057.4]
  assign _T_596 = io_rw_addr == 12'hb18; // @[CSR.scala 177:73:@3058.4]
  assign _T_598 = io_rw_addr == 12'hb98; // @[CSR.scala 177:73:@3059.4]
  assign _T_600 = io_rw_addr == 12'hb19; // @[CSR.scala 177:73:@3060.4]
  assign _T_602 = io_rw_addr == 12'hb99; // @[CSR.scala 177:73:@3061.4]
  assign _T_604 = io_rw_addr == 12'hb1a; // @[CSR.scala 177:73:@3062.4]
  assign _T_606 = io_rw_addr == 12'hb9a; // @[CSR.scala 177:73:@3063.4]
  assign _T_608 = io_rw_addr == 12'hb1b; // @[CSR.scala 177:73:@3064.4]
  assign _T_610 = io_rw_addr == 12'hb9b; // @[CSR.scala 177:73:@3065.4]
  assign _T_612 = io_rw_addr == 12'hb1c; // @[CSR.scala 177:73:@3066.4]
  assign _T_614 = io_rw_addr == 12'hb9c; // @[CSR.scala 177:73:@3067.4]
  assign _T_616 = io_rw_addr == 12'hb1d; // @[CSR.scala 177:73:@3068.4]
  assign _T_618 = io_rw_addr == 12'hb9d; // @[CSR.scala 177:73:@3069.4]
  assign _T_620 = io_rw_addr == 12'hb1e; // @[CSR.scala 177:73:@3070.4]
  assign _T_622 = io_rw_addr == 12'hb9e; // @[CSR.scala 177:73:@3071.4]
  assign _T_624 = io_rw_addr == 12'hb1f; // @[CSR.scala 177:73:@3072.4]
  assign _T_626 = io_rw_addr == 12'hb9f; // @[CSR.scala 177:73:@3073.4]
  assign _T_628 = io_rw_addr == 12'hb20; // @[CSR.scala 177:73:@3074.4]
  assign _T_630 = io_rw_addr == 12'hba0; // @[CSR.scala 177:73:@3075.4]
  assign _T_632 = io_rw_addr == 12'hb21; // @[CSR.scala 177:73:@3076.4]
  assign _T_634 = io_rw_addr == 12'hba1; // @[CSR.scala 177:73:@3077.4]
  assign _T_636 = io_rw_addr == 12'hb22; // @[CSR.scala 177:73:@3078.4]
  assign _T_638 = io_rw_addr == 12'hba2; // @[CSR.scala 177:73:@3079.4]
  assign _T_640 = io_rw_addr == 12'hb80; // @[CSR.scala 177:73:@3080.4]
  assign _T_642 = io_rw_addr == 12'hb82; // @[CSR.scala 177:73:@3081.4]
  assign _T_643 = io_rw_addr[9:8]; // @[CSR.scala 179:54:@3082.4]
  assign priv_sufficient = reg_mstatus_prv >= _T_643; // @[CSR.scala 179:41:@3083.4]
  assign _T_644 = io_rw_addr[11:10]; // @[CSR.scala 180:29:@3084.4]
  assign _T_645 = ~ _T_644; // @[CSR.scala 180:37:@3085.4]
  assign read_only = _T_645 == 2'h0; // @[CSR.scala 180:37:@3086.4]
  assign _T_647 = io_rw_cmd != 3'h5; // @[CSR.scala 181:38:@3087.4]
  assign _T_648 = cpu_ren & _T_647; // @[CSR.scala 181:25:@3088.4]
  assign cpu_wen = _T_648 & priv_sufficient; // @[CSR.scala 181:48:@3089.4]
  assign _T_650 = read_only == 1'h0; // @[CSR.scala 182:24:@3090.4]
  assign wen = cpu_wen & _T_650; // @[CSR.scala 182:21:@3091.4]
  assign _T_651 = io_rw_cmd == 3'h2; // @[Util.scala 23:47:@3092.4]
  assign _T_652 = io_rw_cmd == 3'h3; // @[Util.scala 23:47:@3093.4]
  assign _T_653 = _T_651 | _T_652; // @[Util.scala 23:62:@3094.4]
  assign _T_655 = _T_653 ? io_rw_rdata : 32'h0; // @[CSR.scala 281:9:@3095.4]
  assign _T_656 = _T_655 | io_rw_wdata; // @[CSR.scala 281:49:@3096.4]
  assign _T_659 = _T_652 ? io_rw_wdata : 32'h0; // @[CSR.scala 281:64:@3098.4]
  assign _T_660 = ~ _T_659; // @[CSR.scala 281:60:@3099.4]
  assign wdata = _T_656 & _T_660; // @[CSR.scala 281:58:@3100.4]
  assign _T_662 = io_rw_addr[2:0]; // @[CSR.scala 185:33:@3101.4]
  assign opcode = 8'h1 << _T_662; // @[CSR.scala 185:20:@3102.4]
  assign _T_663 = opcode[0]; // @[CSR.scala 186:40:@3103.4]
  assign insn_call = system_insn & _T_663; // @[CSR.scala 186:31:@3104.4]
  assign _T_664 = opcode[1]; // @[CSR.scala 187:41:@3105.4]
  assign insn_break = system_insn & _T_664; // @[CSR.scala 187:32:@3106.4]
  assign _T_665 = opcode[2]; // @[CSR.scala 188:39:@3107.4]
  assign _T_666 = system_insn & _T_665; // @[CSR.scala 188:30:@3108.4]
  assign insn_ret = _T_666 & priv_sufficient; // @[CSR.scala 188:43:@3109.4]
  assign _T_940 = insn_call | insn_break; // @[CSR.scala 199:24:@3308.4]
  assign _T_942 = {{1'd0}, insn_ret}; // @[Bitwise.scala 48:55:@3311.4]
  assign _T_944 = _T_942 <= 2'h1; // @[CSR.scala 201:50:@3312.4]
  assign _T_946 = _T_944 | reset; // @[CSR.scala 201:9:@3314.4]
  assign _T_948 = _T_946 == 1'h0; // @[CSR.scala 201:9:@3315.4]
  assign _T_951 = io_rw_addr[10]; // @[CSR.scala 208:32:@3324.4]
  assign _T_953 = _T_951 == 1'h0; // @[CSR.scala 208:21:@3325.4]
  assign _T_954 = insn_ret & _T_953; // @[CSR.scala 208:18:@3326.4]
  assign _GEN_3 = _T_954 ? reg_mstatus_mpie : reg_mstatus_mie; // @[CSR.scala 208:38:@3327.4]
  assign _GEN_4 = _T_954 ? 1'h1 : reg_mstatus_mpie; // @[CSR.scala 208:38:@3327.4]
  assign new_prv = _T_954 ? 2'h3 : reg_mstatus_prv; // @[CSR.scala 208:38:@3327.4]
  assign _GEN_148 = {{2'd0}, reg_mstatus_prv}; // @[CSR.scala 218:35:@3335.6]
  assign _T_958 = _GEN_148 + 4'h8; // @[CSR.scala 218:35:@3335.6]
  assign _T_959 = _GEN_148 + 4'h8; // @[CSR.scala 218:35:@3336.6]
  assign _GEN_7 = insn_call ? 32'h80000004 : reg_mepc; // @[CSR.scala 216:18:@3333.4]
  assign _GEN_8 = insn_call ? {{28'd0}, _T_959} : reg_mcause; // @[CSR.scala 216:18:@3333.4]
  assign _GEN_9 = insn_call ? io_pc : reg_mepc; // @[CSR.scala 216:18:@3333.4]
  assign _GEN_10 = insn_break ? 32'h80000004 : _GEN_7; // @[CSR.scala 223:19:@3340.4]
  assign _GEN_11 = insn_break ? 32'h3 : _GEN_8; // @[CSR.scala 223:19:@3340.4]
  assign _GEN_12 = insn_break ? io_pc : _GEN_9; // @[CSR.scala 223:19:@3340.4]
  assign _GEN_14 = io_xcpt ? io_cause : _GEN_11; // @[CSR.scala 229:17:@3345.4]
  assign _GEN_15 = io_xcpt ? io_pc : _GEN_12; // @[CSR.scala 229:17:@3345.4]
  assign _GEN_16 = io_xcpt ? io_tval : reg_mtval; // @[CSR.scala 229:17:@3345.4]
  assign _T_965 = _T_478 ? _T_249 : 64'h0; // @[Mux.scala 19:72:@3353.4]
  assign _T_967 = _T_480 ? _T_261 : 64'h0; // @[Mux.scala 19:72:@3354.4]
  assign _T_969 = _T_482 ? 16'h8000 : 16'h0; // @[Mux.scala 19:72:@3355.4]
  assign _T_975 = _T_488 ? 31'h40000100 : 31'h0; // @[Mux.scala 19:72:@3358.4]
  assign _T_977 = _T_490 ? read_mstatus : 32'h0; // @[Mux.scala 19:72:@3359.4]
  assign _T_979 = _T_492 ? 9'h100 : 9'h0; // @[Mux.scala 19:72:@3360.4]
  assign _T_981 = _T_494 ? _T_468 : 16'h0; // @[Mux.scala 19:72:@3361.4]
  assign _T_983 = _T_496 ? _T_474 : 16'h0; // @[Mux.scala 19:72:@3362.4]
  assign _T_985 = _T_498 ? reg_mscratch : 32'h0; // @[Mux.scala 19:72:@3363.4]
  assign _T_987 = _T_500 ? reg_mepc : 32'h0; // @[Mux.scala 19:72:@3364.4]
  assign _T_989 = _T_502 ? reg_mtval : 32'h0; // @[Mux.scala 19:72:@3365.4]
  assign _T_991 = _T_504 ? reg_mcause : 32'h0; // @[Mux.scala 19:72:@3366.4]
  assign _T_995 = _T_508 ? reg_dscratch : 32'h0; // @[Mux.scala 19:72:@3368.4]
  assign _T_997 = _T_510 ? reg_medeleg : 32'h0; // @[Mux.scala 19:72:@3369.4]
  assign _T_999 = _T_512 ? _T_264 : 40'h0; // @[Mux.scala 19:72:@3370.4]
  assign _T_1001 = _T_514 ? _T_264 : 40'h0; // @[Mux.scala 19:72:@3371.4]
  assign _T_1003 = _T_516 ? _T_267 : 40'h0; // @[Mux.scala 19:72:@3372.4]
  assign _T_1005 = _T_518 ? _T_267 : 40'h0; // @[Mux.scala 19:72:@3373.4]
  assign _T_1007 = _T_520 ? _T_270 : 40'h0; // @[Mux.scala 19:72:@3374.4]
  assign _T_1009 = _T_522 ? _T_270 : 40'h0; // @[Mux.scala 19:72:@3375.4]
  assign _T_1011 = _T_524 ? _T_273 : 40'h0; // @[Mux.scala 19:72:@3376.4]
  assign _T_1013 = _T_526 ? _T_273 : 40'h0; // @[Mux.scala 19:72:@3377.4]
  assign _T_1015 = _T_528 ? _T_276 : 40'h0; // @[Mux.scala 19:72:@3378.4]
  assign _T_1017 = _T_530 ? _T_276 : 40'h0; // @[Mux.scala 19:72:@3379.4]
  assign _T_1019 = _T_532 ? _T_279 : 40'h0; // @[Mux.scala 19:72:@3380.4]
  assign _T_1021 = _T_534 ? _T_279 : 40'h0; // @[Mux.scala 19:72:@3381.4]
  assign _T_1023 = _T_536 ? _T_282 : 40'h0; // @[Mux.scala 19:72:@3382.4]
  assign _T_1025 = _T_538 ? _T_282 : 40'h0; // @[Mux.scala 19:72:@3383.4]
  assign _T_1027 = _T_540 ? _T_285 : 40'h0; // @[Mux.scala 19:72:@3384.4]
  assign _T_1029 = _T_542 ? _T_285 : 40'h0; // @[Mux.scala 19:72:@3385.4]
  assign _T_1031 = _T_544 ? _T_288 : 40'h0; // @[Mux.scala 19:72:@3386.4]
  assign _T_1033 = _T_546 ? _T_288 : 40'h0; // @[Mux.scala 19:72:@3387.4]
  assign _T_1035 = _T_548 ? _T_291 : 40'h0; // @[Mux.scala 19:72:@3388.4]
  assign _T_1037 = _T_550 ? _T_291 : 40'h0; // @[Mux.scala 19:72:@3389.4]
  assign _T_1039 = _T_552 ? _T_294 : 40'h0; // @[Mux.scala 19:72:@3390.4]
  assign _T_1041 = _T_554 ? _T_294 : 40'h0; // @[Mux.scala 19:72:@3391.4]
  assign _T_1043 = _T_556 ? _T_297 : 40'h0; // @[Mux.scala 19:72:@3392.4]
  assign _T_1045 = _T_558 ? _T_297 : 40'h0; // @[Mux.scala 19:72:@3393.4]
  assign _T_1047 = _T_560 ? _T_300 : 40'h0; // @[Mux.scala 19:72:@3394.4]
  assign _T_1049 = _T_562 ? _T_300 : 40'h0; // @[Mux.scala 19:72:@3395.4]
  assign _T_1051 = _T_564 ? _T_303 : 40'h0; // @[Mux.scala 19:72:@3396.4]
  assign _T_1053 = _T_566 ? _T_303 : 40'h0; // @[Mux.scala 19:72:@3397.4]
  assign _T_1055 = _T_568 ? _T_306 : 40'h0; // @[Mux.scala 19:72:@3398.4]
  assign _T_1057 = _T_570 ? _T_306 : 40'h0; // @[Mux.scala 19:72:@3399.4]
  assign _T_1059 = _T_572 ? _T_309 : 40'h0; // @[Mux.scala 19:72:@3400.4]
  assign _T_1061 = _T_574 ? _T_309 : 40'h0; // @[Mux.scala 19:72:@3401.4]
  assign _T_1063 = _T_576 ? _T_312 : 40'h0; // @[Mux.scala 19:72:@3402.4]
  assign _T_1065 = _T_578 ? _T_312 : 40'h0; // @[Mux.scala 19:72:@3403.4]
  assign _T_1067 = _T_580 ? _T_315 : 40'h0; // @[Mux.scala 19:72:@3404.4]
  assign _T_1069 = _T_582 ? _T_315 : 40'h0; // @[Mux.scala 19:72:@3405.4]
  assign _T_1071 = _T_584 ? _T_318 : 40'h0; // @[Mux.scala 19:72:@3406.4]
  assign _T_1073 = _T_586 ? _T_318 : 40'h0; // @[Mux.scala 19:72:@3407.4]
  assign _T_1075 = _T_588 ? _T_321 : 40'h0; // @[Mux.scala 19:72:@3408.4]
  assign _T_1077 = _T_590 ? _T_321 : 40'h0; // @[Mux.scala 19:72:@3409.4]
  assign _T_1079 = _T_592 ? _T_324 : 40'h0; // @[Mux.scala 19:72:@3410.4]
  assign _T_1081 = _T_594 ? _T_324 : 40'h0; // @[Mux.scala 19:72:@3411.4]
  assign _T_1083 = _T_596 ? _T_327 : 40'h0; // @[Mux.scala 19:72:@3412.4]
  assign _T_1085 = _T_598 ? _T_327 : 40'h0; // @[Mux.scala 19:72:@3413.4]
  assign _T_1087 = _T_600 ? _T_330 : 40'h0; // @[Mux.scala 19:72:@3414.4]
  assign _T_1089 = _T_602 ? _T_330 : 40'h0; // @[Mux.scala 19:72:@3415.4]
  assign _T_1091 = _T_604 ? _T_333 : 40'h0; // @[Mux.scala 19:72:@3416.4]
  assign _T_1093 = _T_606 ? _T_333 : 40'h0; // @[Mux.scala 19:72:@3417.4]
  assign _T_1095 = _T_608 ? _T_336 : 40'h0; // @[Mux.scala 19:72:@3418.4]
  assign _T_1097 = _T_610 ? _T_336 : 40'h0; // @[Mux.scala 19:72:@3419.4]
  assign _T_1099 = _T_612 ? _T_339 : 40'h0; // @[Mux.scala 19:72:@3420.4]
  assign _T_1101 = _T_614 ? _T_339 : 40'h0; // @[Mux.scala 19:72:@3421.4]
  assign _T_1103 = _T_616 ? _T_342 : 40'h0; // @[Mux.scala 19:72:@3422.4]
  assign _T_1105 = _T_618 ? _T_342 : 40'h0; // @[Mux.scala 19:72:@3423.4]
  assign _T_1107 = _T_620 ? _T_345 : 40'h0; // @[Mux.scala 19:72:@3424.4]
  assign _T_1109 = _T_622 ? _T_345 : 40'h0; // @[Mux.scala 19:72:@3425.4]
  assign _T_1111 = _T_624 ? _T_348 : 40'h0; // @[Mux.scala 19:72:@3426.4]
  assign _T_1113 = _T_626 ? _T_348 : 40'h0; // @[Mux.scala 19:72:@3427.4]
  assign _T_1115 = _T_628 ? _T_351 : 40'h0; // @[Mux.scala 19:72:@3428.4]
  assign _T_1117 = _T_630 ? _T_351 : 40'h0; // @[Mux.scala 19:72:@3429.4]
  assign _T_1119 = _T_632 ? _T_354 : 40'h0; // @[Mux.scala 19:72:@3430.4]
  assign _T_1121 = _T_634 ? _T_354 : 40'h0; // @[Mux.scala 19:72:@3431.4]
  assign _T_1123 = _T_636 ? _T_357 : 40'h0; // @[Mux.scala 19:72:@3432.4]
  assign _T_1125 = _T_638 ? _T_357 : 40'h0; // @[Mux.scala 19:72:@3433.4]
  assign _T_1130 = _T_965 | _T_967; // @[Mux.scala 19:72:@3436.4]
  assign _GEN_149 = {{48'd0}, _T_969}; // @[Mux.scala 19:72:@3437.4]
  assign _T_1131 = _T_1130 | _GEN_149; // @[Mux.scala 19:72:@3437.4]
  assign _GEN_150 = {{33'd0}, _T_975}; // @[Mux.scala 19:72:@3440.4]
  assign _T_1134 = _T_1131 | _GEN_150; // @[Mux.scala 19:72:@3440.4]
  assign _GEN_151 = {{32'd0}, _T_977}; // @[Mux.scala 19:72:@3441.4]
  assign _T_1135 = _T_1134 | _GEN_151; // @[Mux.scala 19:72:@3441.4]
  assign _GEN_152 = {{55'd0}, _T_979}; // @[Mux.scala 19:72:@3442.4]
  assign _T_1136 = _T_1135 | _GEN_152; // @[Mux.scala 19:72:@3442.4]
  assign _GEN_153 = {{48'd0}, _T_981}; // @[Mux.scala 19:72:@3443.4]
  assign _T_1137 = _T_1136 | _GEN_153; // @[Mux.scala 19:72:@3443.4]
  assign _GEN_154 = {{48'd0}, _T_983}; // @[Mux.scala 19:72:@3444.4]
  assign _T_1138 = _T_1137 | _GEN_154; // @[Mux.scala 19:72:@3444.4]
  assign _GEN_155 = {{32'd0}, _T_985}; // @[Mux.scala 19:72:@3445.4]
  assign _T_1139 = _T_1138 | _GEN_155; // @[Mux.scala 19:72:@3445.4]
  assign _GEN_156 = {{32'd0}, _T_987}; // @[Mux.scala 19:72:@3446.4]
  assign _T_1140 = _T_1139 | _GEN_156; // @[Mux.scala 19:72:@3446.4]
  assign _GEN_157 = {{32'd0}, _T_989}; // @[Mux.scala 19:72:@3447.4]
  assign _T_1141 = _T_1140 | _GEN_157; // @[Mux.scala 19:72:@3447.4]
  assign _GEN_158 = {{32'd0}, _T_991}; // @[Mux.scala 19:72:@3448.4]
  assign _T_1142 = _T_1141 | _GEN_158; // @[Mux.scala 19:72:@3448.4]
  assign _GEN_159 = {{32'd0}, _T_995}; // @[Mux.scala 19:72:@3450.4]
  assign _T_1144 = _T_1142 | _GEN_159; // @[Mux.scala 19:72:@3450.4]
  assign _GEN_160 = {{32'd0}, _T_997}; // @[Mux.scala 19:72:@3451.4]
  assign _T_1145 = _T_1144 | _GEN_160; // @[Mux.scala 19:72:@3451.4]
  assign _GEN_161 = {{24'd0}, _T_999}; // @[Mux.scala 19:72:@3452.4]
  assign _T_1146 = _T_1145 | _GEN_161; // @[Mux.scala 19:72:@3452.4]
  assign _GEN_162 = {{24'd0}, _T_1001}; // @[Mux.scala 19:72:@3453.4]
  assign _T_1147 = _T_1146 | _GEN_162; // @[Mux.scala 19:72:@3453.4]
  assign _GEN_163 = {{24'd0}, _T_1003}; // @[Mux.scala 19:72:@3454.4]
  assign _T_1148 = _T_1147 | _GEN_163; // @[Mux.scala 19:72:@3454.4]
  assign _GEN_164 = {{24'd0}, _T_1005}; // @[Mux.scala 19:72:@3455.4]
  assign _T_1149 = _T_1148 | _GEN_164; // @[Mux.scala 19:72:@3455.4]
  assign _GEN_165 = {{24'd0}, _T_1007}; // @[Mux.scala 19:72:@3456.4]
  assign _T_1150 = _T_1149 | _GEN_165; // @[Mux.scala 19:72:@3456.4]
  assign _GEN_166 = {{24'd0}, _T_1009}; // @[Mux.scala 19:72:@3457.4]
  assign _T_1151 = _T_1150 | _GEN_166; // @[Mux.scala 19:72:@3457.4]
  assign _GEN_167 = {{24'd0}, _T_1011}; // @[Mux.scala 19:72:@3458.4]
  assign _T_1152 = _T_1151 | _GEN_167; // @[Mux.scala 19:72:@3458.4]
  assign _GEN_168 = {{24'd0}, _T_1013}; // @[Mux.scala 19:72:@3459.4]
  assign _T_1153 = _T_1152 | _GEN_168; // @[Mux.scala 19:72:@3459.4]
  assign _GEN_169 = {{24'd0}, _T_1015}; // @[Mux.scala 19:72:@3460.4]
  assign _T_1154 = _T_1153 | _GEN_169; // @[Mux.scala 19:72:@3460.4]
  assign _GEN_170 = {{24'd0}, _T_1017}; // @[Mux.scala 19:72:@3461.4]
  assign _T_1155 = _T_1154 | _GEN_170; // @[Mux.scala 19:72:@3461.4]
  assign _GEN_171 = {{24'd0}, _T_1019}; // @[Mux.scala 19:72:@3462.4]
  assign _T_1156 = _T_1155 | _GEN_171; // @[Mux.scala 19:72:@3462.4]
  assign _GEN_172 = {{24'd0}, _T_1021}; // @[Mux.scala 19:72:@3463.4]
  assign _T_1157 = _T_1156 | _GEN_172; // @[Mux.scala 19:72:@3463.4]
  assign _GEN_173 = {{24'd0}, _T_1023}; // @[Mux.scala 19:72:@3464.4]
  assign _T_1158 = _T_1157 | _GEN_173; // @[Mux.scala 19:72:@3464.4]
  assign _GEN_174 = {{24'd0}, _T_1025}; // @[Mux.scala 19:72:@3465.4]
  assign _T_1159 = _T_1158 | _GEN_174; // @[Mux.scala 19:72:@3465.4]
  assign _GEN_175 = {{24'd0}, _T_1027}; // @[Mux.scala 19:72:@3466.4]
  assign _T_1160 = _T_1159 | _GEN_175; // @[Mux.scala 19:72:@3466.4]
  assign _GEN_176 = {{24'd0}, _T_1029}; // @[Mux.scala 19:72:@3467.4]
  assign _T_1161 = _T_1160 | _GEN_176; // @[Mux.scala 19:72:@3467.4]
  assign _GEN_177 = {{24'd0}, _T_1031}; // @[Mux.scala 19:72:@3468.4]
  assign _T_1162 = _T_1161 | _GEN_177; // @[Mux.scala 19:72:@3468.4]
  assign _GEN_178 = {{24'd0}, _T_1033}; // @[Mux.scala 19:72:@3469.4]
  assign _T_1163 = _T_1162 | _GEN_178; // @[Mux.scala 19:72:@3469.4]
  assign _GEN_179 = {{24'd0}, _T_1035}; // @[Mux.scala 19:72:@3470.4]
  assign _T_1164 = _T_1163 | _GEN_179; // @[Mux.scala 19:72:@3470.4]
  assign _GEN_180 = {{24'd0}, _T_1037}; // @[Mux.scala 19:72:@3471.4]
  assign _T_1165 = _T_1164 | _GEN_180; // @[Mux.scala 19:72:@3471.4]
  assign _GEN_181 = {{24'd0}, _T_1039}; // @[Mux.scala 19:72:@3472.4]
  assign _T_1166 = _T_1165 | _GEN_181; // @[Mux.scala 19:72:@3472.4]
  assign _GEN_182 = {{24'd0}, _T_1041}; // @[Mux.scala 19:72:@3473.4]
  assign _T_1167 = _T_1166 | _GEN_182; // @[Mux.scala 19:72:@3473.4]
  assign _GEN_183 = {{24'd0}, _T_1043}; // @[Mux.scala 19:72:@3474.4]
  assign _T_1168 = _T_1167 | _GEN_183; // @[Mux.scala 19:72:@3474.4]
  assign _GEN_184 = {{24'd0}, _T_1045}; // @[Mux.scala 19:72:@3475.4]
  assign _T_1169 = _T_1168 | _GEN_184; // @[Mux.scala 19:72:@3475.4]
  assign _GEN_185 = {{24'd0}, _T_1047}; // @[Mux.scala 19:72:@3476.4]
  assign _T_1170 = _T_1169 | _GEN_185; // @[Mux.scala 19:72:@3476.4]
  assign _GEN_186 = {{24'd0}, _T_1049}; // @[Mux.scala 19:72:@3477.4]
  assign _T_1171 = _T_1170 | _GEN_186; // @[Mux.scala 19:72:@3477.4]
  assign _GEN_187 = {{24'd0}, _T_1051}; // @[Mux.scala 19:72:@3478.4]
  assign _T_1172 = _T_1171 | _GEN_187; // @[Mux.scala 19:72:@3478.4]
  assign _GEN_188 = {{24'd0}, _T_1053}; // @[Mux.scala 19:72:@3479.4]
  assign _T_1173 = _T_1172 | _GEN_188; // @[Mux.scala 19:72:@3479.4]
  assign _GEN_189 = {{24'd0}, _T_1055}; // @[Mux.scala 19:72:@3480.4]
  assign _T_1174 = _T_1173 | _GEN_189; // @[Mux.scala 19:72:@3480.4]
  assign _GEN_190 = {{24'd0}, _T_1057}; // @[Mux.scala 19:72:@3481.4]
  assign _T_1175 = _T_1174 | _GEN_190; // @[Mux.scala 19:72:@3481.4]
  assign _GEN_191 = {{24'd0}, _T_1059}; // @[Mux.scala 19:72:@3482.4]
  assign _T_1176 = _T_1175 | _GEN_191; // @[Mux.scala 19:72:@3482.4]
  assign _GEN_192 = {{24'd0}, _T_1061}; // @[Mux.scala 19:72:@3483.4]
  assign _T_1177 = _T_1176 | _GEN_192; // @[Mux.scala 19:72:@3483.4]
  assign _GEN_193 = {{24'd0}, _T_1063}; // @[Mux.scala 19:72:@3484.4]
  assign _T_1178 = _T_1177 | _GEN_193; // @[Mux.scala 19:72:@3484.4]
  assign _GEN_194 = {{24'd0}, _T_1065}; // @[Mux.scala 19:72:@3485.4]
  assign _T_1179 = _T_1178 | _GEN_194; // @[Mux.scala 19:72:@3485.4]
  assign _GEN_195 = {{24'd0}, _T_1067}; // @[Mux.scala 19:72:@3486.4]
  assign _T_1180 = _T_1179 | _GEN_195; // @[Mux.scala 19:72:@3486.4]
  assign _GEN_196 = {{24'd0}, _T_1069}; // @[Mux.scala 19:72:@3487.4]
  assign _T_1181 = _T_1180 | _GEN_196; // @[Mux.scala 19:72:@3487.4]
  assign _GEN_197 = {{24'd0}, _T_1071}; // @[Mux.scala 19:72:@3488.4]
  assign _T_1182 = _T_1181 | _GEN_197; // @[Mux.scala 19:72:@3488.4]
  assign _GEN_198 = {{24'd0}, _T_1073}; // @[Mux.scala 19:72:@3489.4]
  assign _T_1183 = _T_1182 | _GEN_198; // @[Mux.scala 19:72:@3489.4]
  assign _GEN_199 = {{24'd0}, _T_1075}; // @[Mux.scala 19:72:@3490.4]
  assign _T_1184 = _T_1183 | _GEN_199; // @[Mux.scala 19:72:@3490.4]
  assign _GEN_200 = {{24'd0}, _T_1077}; // @[Mux.scala 19:72:@3491.4]
  assign _T_1185 = _T_1184 | _GEN_200; // @[Mux.scala 19:72:@3491.4]
  assign _GEN_201 = {{24'd0}, _T_1079}; // @[Mux.scala 19:72:@3492.4]
  assign _T_1186 = _T_1185 | _GEN_201; // @[Mux.scala 19:72:@3492.4]
  assign _GEN_202 = {{24'd0}, _T_1081}; // @[Mux.scala 19:72:@3493.4]
  assign _T_1187 = _T_1186 | _GEN_202; // @[Mux.scala 19:72:@3493.4]
  assign _GEN_203 = {{24'd0}, _T_1083}; // @[Mux.scala 19:72:@3494.4]
  assign _T_1188 = _T_1187 | _GEN_203; // @[Mux.scala 19:72:@3494.4]
  assign _GEN_204 = {{24'd0}, _T_1085}; // @[Mux.scala 19:72:@3495.4]
  assign _T_1189 = _T_1188 | _GEN_204; // @[Mux.scala 19:72:@3495.4]
  assign _GEN_205 = {{24'd0}, _T_1087}; // @[Mux.scala 19:72:@3496.4]
  assign _T_1190 = _T_1189 | _GEN_205; // @[Mux.scala 19:72:@3496.4]
  assign _GEN_206 = {{24'd0}, _T_1089}; // @[Mux.scala 19:72:@3497.4]
  assign _T_1191 = _T_1190 | _GEN_206; // @[Mux.scala 19:72:@3497.4]
  assign _GEN_207 = {{24'd0}, _T_1091}; // @[Mux.scala 19:72:@3498.4]
  assign _T_1192 = _T_1191 | _GEN_207; // @[Mux.scala 19:72:@3498.4]
  assign _GEN_208 = {{24'd0}, _T_1093}; // @[Mux.scala 19:72:@3499.4]
  assign _T_1193 = _T_1192 | _GEN_208; // @[Mux.scala 19:72:@3499.4]
  assign _GEN_209 = {{24'd0}, _T_1095}; // @[Mux.scala 19:72:@3500.4]
  assign _T_1194 = _T_1193 | _GEN_209; // @[Mux.scala 19:72:@3500.4]
  assign _GEN_210 = {{24'd0}, _T_1097}; // @[Mux.scala 19:72:@3501.4]
  assign _T_1195 = _T_1194 | _GEN_210; // @[Mux.scala 19:72:@3501.4]
  assign _GEN_211 = {{24'd0}, _T_1099}; // @[Mux.scala 19:72:@3502.4]
  assign _T_1196 = _T_1195 | _GEN_211; // @[Mux.scala 19:72:@3502.4]
  assign _GEN_212 = {{24'd0}, _T_1101}; // @[Mux.scala 19:72:@3503.4]
  assign _T_1197 = _T_1196 | _GEN_212; // @[Mux.scala 19:72:@3503.4]
  assign _GEN_213 = {{24'd0}, _T_1103}; // @[Mux.scala 19:72:@3504.4]
  assign _T_1198 = _T_1197 | _GEN_213; // @[Mux.scala 19:72:@3504.4]
  assign _GEN_214 = {{24'd0}, _T_1105}; // @[Mux.scala 19:72:@3505.4]
  assign _T_1199 = _T_1198 | _GEN_214; // @[Mux.scala 19:72:@3505.4]
  assign _GEN_215 = {{24'd0}, _T_1107}; // @[Mux.scala 19:72:@3506.4]
  assign _T_1200 = _T_1199 | _GEN_215; // @[Mux.scala 19:72:@3506.4]
  assign _GEN_216 = {{24'd0}, _T_1109}; // @[Mux.scala 19:72:@3507.4]
  assign _T_1201 = _T_1200 | _GEN_216; // @[Mux.scala 19:72:@3507.4]
  assign _GEN_217 = {{24'd0}, _T_1111}; // @[Mux.scala 19:72:@3508.4]
  assign _T_1202 = _T_1201 | _GEN_217; // @[Mux.scala 19:72:@3508.4]
  assign _GEN_218 = {{24'd0}, _T_1113}; // @[Mux.scala 19:72:@3509.4]
  assign _T_1203 = _T_1202 | _GEN_218; // @[Mux.scala 19:72:@3509.4]
  assign _GEN_219 = {{24'd0}, _T_1115}; // @[Mux.scala 19:72:@3510.4]
  assign _T_1204 = _T_1203 | _GEN_219; // @[Mux.scala 19:72:@3510.4]
  assign _GEN_220 = {{24'd0}, _T_1117}; // @[Mux.scala 19:72:@3511.4]
  assign _T_1205 = _T_1204 | _GEN_220; // @[Mux.scala 19:72:@3511.4]
  assign _GEN_221 = {{24'd0}, _T_1119}; // @[Mux.scala 19:72:@3512.4]
  assign _T_1206 = _T_1205 | _GEN_221; // @[Mux.scala 19:72:@3512.4]
  assign _GEN_222 = {{24'd0}, _T_1121}; // @[Mux.scala 19:72:@3513.4]
  assign _T_1207 = _T_1206 | _GEN_222; // @[Mux.scala 19:72:@3513.4]
  assign _GEN_223 = {{24'd0}, _T_1123}; // @[Mux.scala 19:72:@3514.4]
  assign _T_1208 = _T_1207 | _GEN_223; // @[Mux.scala 19:72:@3514.4]
  assign _GEN_224 = {{24'd0}, _T_1125}; // @[Mux.scala 19:72:@3515.4]
  assign _T_1209 = _T_1208 | _GEN_224; // @[Mux.scala 19:72:@3515.4]
  assign _T_1220 = wdata[3]; // @[CSR.scala 245:39:@3528.8]
  assign _T_1222 = wdata[7]; // @[CSR.scala 245:39:@3532.8]
  assign _GEN_17 = _T_490 ? _T_1220 : _GEN_3; // @[CSR.scala 244:39:@3522.6]
  assign _GEN_18 = _T_490 ? _T_1222 : _GEN_4; // @[CSR.scala 244:39:@3522.6]
  assign _T_1233 = wdata[15:0]; // @[:@3551.8 :@3552.8]
  assign _T_1235 = _T_1233[3]; // @[CSR.scala 250:35:@3555.8]
  assign _T_1237 = _T_1233[7]; // @[CSR.scala 250:35:@3559.8]
  assign _GEN_19 = _T_494 ? _T_1235 : reg_mip_msip; // @[CSR.scala 249:35:@3549.6]
  assign _GEN_20 = _T_496 ? _T_1235 : reg_mie_msip; // @[CSR.scala 253:35:@3569.6]
  assign _GEN_21 = _T_496 ? _T_1237 : reg_mie_mtip; // @[CSR.scala 253:35:@3569.6]
  assign _T_1253 = wdata[7:0]; // @[CSR.scala 277:47:@3591.8]
  assign _T_1254 = _T_264[31:0]; // @[CSR.scala 277:72:@3592.8]
  assign _T_1255 = {_T_1253,_T_1254}; // @[Cat.scala 30:58:@3593.8]
  assign _GEN_22 = _T_514 ? {{1'd0}, _T_1255} : _T_265; // @[CSR.scala 277:29:@3590.6]
  assign _T_1256 = _T_264[39:32]; // @[CSR.scala 278:45:@3597.8]
  assign _T_1257 = {_T_1256,wdata}; // @[Cat.scala 30:58:@3598.8]
  assign _GEN_23 = _T_512 ? {{1'd0}, _T_1257} : _GEN_22; // @[CSR.scala 278:29:@3596.6]
  assign _T_1259 = _T_267[31:0]; // @[CSR.scala 277:72:@3603.8]
  assign _T_1260 = {_T_1253,_T_1259}; // @[Cat.scala 30:58:@3604.8]
  assign _GEN_24 = _T_518 ? {{1'd0}, _T_1260} : _T_268; // @[CSR.scala 277:29:@3601.6]
  assign _T_1261 = _T_267[39:32]; // @[CSR.scala 278:45:@3608.8]
  assign _T_1262 = {_T_1261,wdata}; // @[Cat.scala 30:58:@3609.8]
  assign _GEN_25 = _T_516 ? {{1'd0}, _T_1262} : _GEN_24; // @[CSR.scala 278:29:@3607.6]
  assign _T_1264 = _T_270[31:0]; // @[CSR.scala 277:72:@3614.8]
  assign _T_1265 = {_T_1253,_T_1264}; // @[Cat.scala 30:58:@3615.8]
  assign _GEN_26 = _T_522 ? {{1'd0}, _T_1265} : _T_271; // @[CSR.scala 277:29:@3612.6]
  assign _T_1266 = _T_270[39:32]; // @[CSR.scala 278:45:@3619.8]
  assign _T_1267 = {_T_1266,wdata}; // @[Cat.scala 30:58:@3620.8]
  assign _GEN_27 = _T_520 ? {{1'd0}, _T_1267} : _GEN_26; // @[CSR.scala 278:29:@3618.6]
  assign _T_1269 = _T_273[31:0]; // @[CSR.scala 277:72:@3625.8]
  assign _T_1270 = {_T_1253,_T_1269}; // @[Cat.scala 30:58:@3626.8]
  assign _GEN_28 = _T_526 ? {{1'd0}, _T_1270} : _T_274; // @[CSR.scala 277:29:@3623.6]
  assign _T_1271 = _T_273[39:32]; // @[CSR.scala 278:45:@3630.8]
  assign _T_1272 = {_T_1271,wdata}; // @[Cat.scala 30:58:@3631.8]
  assign _GEN_29 = _T_524 ? {{1'd0}, _T_1272} : _GEN_28; // @[CSR.scala 278:29:@3629.6]
  assign _T_1274 = _T_276[31:0]; // @[CSR.scala 277:72:@3636.8]
  assign _T_1275 = {_T_1253,_T_1274}; // @[Cat.scala 30:58:@3637.8]
  assign _GEN_30 = _T_530 ? {{1'd0}, _T_1275} : _T_277; // @[CSR.scala 277:29:@3634.6]
  assign _T_1276 = _T_276[39:32]; // @[CSR.scala 278:45:@3641.8]
  assign _T_1277 = {_T_1276,wdata}; // @[Cat.scala 30:58:@3642.8]
  assign _GEN_31 = _T_528 ? {{1'd0}, _T_1277} : _GEN_30; // @[CSR.scala 278:29:@3640.6]
  assign _T_1279 = _T_279[31:0]; // @[CSR.scala 277:72:@3647.8]
  assign _T_1280 = {_T_1253,_T_1279}; // @[Cat.scala 30:58:@3648.8]
  assign _GEN_32 = _T_534 ? {{1'd0}, _T_1280} : _T_280; // @[CSR.scala 277:29:@3645.6]
  assign _T_1281 = _T_279[39:32]; // @[CSR.scala 278:45:@3652.8]
  assign _T_1282 = {_T_1281,wdata}; // @[Cat.scala 30:58:@3653.8]
  assign _GEN_33 = _T_532 ? {{1'd0}, _T_1282} : _GEN_32; // @[CSR.scala 278:29:@3651.6]
  assign _T_1284 = _T_282[31:0]; // @[CSR.scala 277:72:@3658.8]
  assign _T_1285 = {_T_1253,_T_1284}; // @[Cat.scala 30:58:@3659.8]
  assign _GEN_34 = _T_538 ? {{1'd0}, _T_1285} : _T_283; // @[CSR.scala 277:29:@3656.6]
  assign _T_1286 = _T_282[39:32]; // @[CSR.scala 278:45:@3663.8]
  assign _T_1287 = {_T_1286,wdata}; // @[Cat.scala 30:58:@3664.8]
  assign _GEN_35 = _T_536 ? {{1'd0}, _T_1287} : _GEN_34; // @[CSR.scala 278:29:@3662.6]
  assign _T_1289 = _T_285[31:0]; // @[CSR.scala 277:72:@3669.8]
  assign _T_1290 = {_T_1253,_T_1289}; // @[Cat.scala 30:58:@3670.8]
  assign _GEN_36 = _T_542 ? {{1'd0}, _T_1290} : _T_286; // @[CSR.scala 277:29:@3667.6]
  assign _T_1291 = _T_285[39:32]; // @[CSR.scala 278:45:@3674.8]
  assign _T_1292 = {_T_1291,wdata}; // @[Cat.scala 30:58:@3675.8]
  assign _GEN_37 = _T_540 ? {{1'd0}, _T_1292} : _GEN_36; // @[CSR.scala 278:29:@3673.6]
  assign _T_1294 = _T_288[31:0]; // @[CSR.scala 277:72:@3680.8]
  assign _T_1295 = {_T_1253,_T_1294}; // @[Cat.scala 30:58:@3681.8]
  assign _GEN_38 = _T_546 ? {{1'd0}, _T_1295} : _T_289; // @[CSR.scala 277:29:@3678.6]
  assign _T_1296 = _T_288[39:32]; // @[CSR.scala 278:45:@3685.8]
  assign _T_1297 = {_T_1296,wdata}; // @[Cat.scala 30:58:@3686.8]
  assign _GEN_39 = _T_544 ? {{1'd0}, _T_1297} : _GEN_38; // @[CSR.scala 278:29:@3684.6]
  assign _T_1299 = _T_291[31:0]; // @[CSR.scala 277:72:@3691.8]
  assign _T_1300 = {_T_1253,_T_1299}; // @[Cat.scala 30:58:@3692.8]
  assign _GEN_40 = _T_550 ? {{1'd0}, _T_1300} : _T_292; // @[CSR.scala 277:29:@3689.6]
  assign _T_1301 = _T_291[39:32]; // @[CSR.scala 278:45:@3696.8]
  assign _T_1302 = {_T_1301,wdata}; // @[Cat.scala 30:58:@3697.8]
  assign _GEN_41 = _T_548 ? {{1'd0}, _T_1302} : _GEN_40; // @[CSR.scala 278:29:@3695.6]
  assign _T_1304 = _T_294[31:0]; // @[CSR.scala 277:72:@3702.8]
  assign _T_1305 = {_T_1253,_T_1304}; // @[Cat.scala 30:58:@3703.8]
  assign _GEN_42 = _T_554 ? {{1'd0}, _T_1305} : _T_295; // @[CSR.scala 277:29:@3700.6]
  assign _T_1306 = _T_294[39:32]; // @[CSR.scala 278:45:@3707.8]
  assign _T_1307 = {_T_1306,wdata}; // @[Cat.scala 30:58:@3708.8]
  assign _GEN_43 = _T_552 ? {{1'd0}, _T_1307} : _GEN_42; // @[CSR.scala 278:29:@3706.6]
  assign _T_1309 = _T_297[31:0]; // @[CSR.scala 277:72:@3713.8]
  assign _T_1310 = {_T_1253,_T_1309}; // @[Cat.scala 30:58:@3714.8]
  assign _GEN_44 = _T_558 ? {{1'd0}, _T_1310} : _T_298; // @[CSR.scala 277:29:@3711.6]
  assign _T_1311 = _T_297[39:32]; // @[CSR.scala 278:45:@3718.8]
  assign _T_1312 = {_T_1311,wdata}; // @[Cat.scala 30:58:@3719.8]
  assign _GEN_45 = _T_556 ? {{1'd0}, _T_1312} : _GEN_44; // @[CSR.scala 278:29:@3717.6]
  assign _T_1314 = _T_300[31:0]; // @[CSR.scala 277:72:@3724.8]
  assign _T_1315 = {_T_1253,_T_1314}; // @[Cat.scala 30:58:@3725.8]
  assign _GEN_46 = _T_562 ? {{1'd0}, _T_1315} : _T_301; // @[CSR.scala 277:29:@3722.6]
  assign _T_1316 = _T_300[39:32]; // @[CSR.scala 278:45:@3729.8]
  assign _T_1317 = {_T_1316,wdata}; // @[Cat.scala 30:58:@3730.8]
  assign _GEN_47 = _T_560 ? {{1'd0}, _T_1317} : _GEN_46; // @[CSR.scala 278:29:@3728.6]
  assign _T_1319 = _T_303[31:0]; // @[CSR.scala 277:72:@3735.8]
  assign _T_1320 = {_T_1253,_T_1319}; // @[Cat.scala 30:58:@3736.8]
  assign _GEN_48 = _T_566 ? {{1'd0}, _T_1320} : _T_304; // @[CSR.scala 277:29:@3733.6]
  assign _T_1321 = _T_303[39:32]; // @[CSR.scala 278:45:@3740.8]
  assign _T_1322 = {_T_1321,wdata}; // @[Cat.scala 30:58:@3741.8]
  assign _GEN_49 = _T_564 ? {{1'd0}, _T_1322} : _GEN_48; // @[CSR.scala 278:29:@3739.6]
  assign _T_1324 = _T_306[31:0]; // @[CSR.scala 277:72:@3746.8]
  assign _T_1325 = {_T_1253,_T_1324}; // @[Cat.scala 30:58:@3747.8]
  assign _GEN_50 = _T_570 ? {{1'd0}, _T_1325} : _T_307; // @[CSR.scala 277:29:@3744.6]
  assign _T_1326 = _T_306[39:32]; // @[CSR.scala 278:45:@3751.8]
  assign _T_1327 = {_T_1326,wdata}; // @[Cat.scala 30:58:@3752.8]
  assign _GEN_51 = _T_568 ? {{1'd0}, _T_1327} : _GEN_50; // @[CSR.scala 278:29:@3750.6]
  assign _T_1329 = _T_309[31:0]; // @[CSR.scala 277:72:@3757.8]
  assign _T_1330 = {_T_1253,_T_1329}; // @[Cat.scala 30:58:@3758.8]
  assign _GEN_52 = _T_574 ? {{1'd0}, _T_1330} : _T_310; // @[CSR.scala 277:29:@3755.6]
  assign _T_1331 = _T_309[39:32]; // @[CSR.scala 278:45:@3762.8]
  assign _T_1332 = {_T_1331,wdata}; // @[Cat.scala 30:58:@3763.8]
  assign _GEN_53 = _T_572 ? {{1'd0}, _T_1332} : _GEN_52; // @[CSR.scala 278:29:@3761.6]
  assign _T_1334 = _T_312[31:0]; // @[CSR.scala 277:72:@3768.8]
  assign _T_1335 = {_T_1253,_T_1334}; // @[Cat.scala 30:58:@3769.8]
  assign _GEN_54 = _T_578 ? {{1'd0}, _T_1335} : _T_313; // @[CSR.scala 277:29:@3766.6]
  assign _T_1336 = _T_312[39:32]; // @[CSR.scala 278:45:@3773.8]
  assign _T_1337 = {_T_1336,wdata}; // @[Cat.scala 30:58:@3774.8]
  assign _GEN_55 = _T_576 ? {{1'd0}, _T_1337} : _GEN_54; // @[CSR.scala 278:29:@3772.6]
  assign _T_1339 = _T_315[31:0]; // @[CSR.scala 277:72:@3779.8]
  assign _T_1340 = {_T_1253,_T_1339}; // @[Cat.scala 30:58:@3780.8]
  assign _GEN_56 = _T_582 ? {{1'd0}, _T_1340} : _T_316; // @[CSR.scala 277:29:@3777.6]
  assign _T_1341 = _T_315[39:32]; // @[CSR.scala 278:45:@3784.8]
  assign _T_1342 = {_T_1341,wdata}; // @[Cat.scala 30:58:@3785.8]
  assign _GEN_57 = _T_580 ? {{1'd0}, _T_1342} : _GEN_56; // @[CSR.scala 278:29:@3783.6]
  assign _T_1344 = _T_318[31:0]; // @[CSR.scala 277:72:@3790.8]
  assign _T_1345 = {_T_1253,_T_1344}; // @[Cat.scala 30:58:@3791.8]
  assign _GEN_58 = _T_586 ? {{1'd0}, _T_1345} : _T_319; // @[CSR.scala 277:29:@3788.6]
  assign _T_1346 = _T_318[39:32]; // @[CSR.scala 278:45:@3795.8]
  assign _T_1347 = {_T_1346,wdata}; // @[Cat.scala 30:58:@3796.8]
  assign _GEN_59 = _T_584 ? {{1'd0}, _T_1347} : _GEN_58; // @[CSR.scala 278:29:@3794.6]
  assign _T_1349 = _T_321[31:0]; // @[CSR.scala 277:72:@3801.8]
  assign _T_1350 = {_T_1253,_T_1349}; // @[Cat.scala 30:58:@3802.8]
  assign _GEN_60 = _T_590 ? {{1'd0}, _T_1350} : _T_322; // @[CSR.scala 277:29:@3799.6]
  assign _T_1351 = _T_321[39:32]; // @[CSR.scala 278:45:@3806.8]
  assign _T_1352 = {_T_1351,wdata}; // @[Cat.scala 30:58:@3807.8]
  assign _GEN_61 = _T_588 ? {{1'd0}, _T_1352} : _GEN_60; // @[CSR.scala 278:29:@3805.6]
  assign _T_1354 = _T_324[31:0]; // @[CSR.scala 277:72:@3812.8]
  assign _T_1355 = {_T_1253,_T_1354}; // @[Cat.scala 30:58:@3813.8]
  assign _GEN_62 = _T_594 ? {{1'd0}, _T_1355} : _T_325; // @[CSR.scala 277:29:@3810.6]
  assign _T_1356 = _T_324[39:32]; // @[CSR.scala 278:45:@3817.8]
  assign _T_1357 = {_T_1356,wdata}; // @[Cat.scala 30:58:@3818.8]
  assign _GEN_63 = _T_592 ? {{1'd0}, _T_1357} : _GEN_62; // @[CSR.scala 278:29:@3816.6]
  assign _T_1359 = _T_327[31:0]; // @[CSR.scala 277:72:@3823.8]
  assign _T_1360 = {_T_1253,_T_1359}; // @[Cat.scala 30:58:@3824.8]
  assign _GEN_64 = _T_598 ? {{1'd0}, _T_1360} : _T_328; // @[CSR.scala 277:29:@3821.6]
  assign _T_1361 = _T_327[39:32]; // @[CSR.scala 278:45:@3828.8]
  assign _T_1362 = {_T_1361,wdata}; // @[Cat.scala 30:58:@3829.8]
  assign _GEN_65 = _T_596 ? {{1'd0}, _T_1362} : _GEN_64; // @[CSR.scala 278:29:@3827.6]
  assign _T_1364 = _T_330[31:0]; // @[CSR.scala 277:72:@3834.8]
  assign _T_1365 = {_T_1253,_T_1364}; // @[Cat.scala 30:58:@3835.8]
  assign _GEN_66 = _T_602 ? {{1'd0}, _T_1365} : _T_331; // @[CSR.scala 277:29:@3832.6]
  assign _T_1366 = _T_330[39:32]; // @[CSR.scala 278:45:@3839.8]
  assign _T_1367 = {_T_1366,wdata}; // @[Cat.scala 30:58:@3840.8]
  assign _GEN_67 = _T_600 ? {{1'd0}, _T_1367} : _GEN_66; // @[CSR.scala 278:29:@3838.6]
  assign _T_1369 = _T_333[31:0]; // @[CSR.scala 277:72:@3845.8]
  assign _T_1370 = {_T_1253,_T_1369}; // @[Cat.scala 30:58:@3846.8]
  assign _GEN_68 = _T_606 ? {{1'd0}, _T_1370} : _T_334; // @[CSR.scala 277:29:@3843.6]
  assign _T_1371 = _T_333[39:32]; // @[CSR.scala 278:45:@3850.8]
  assign _T_1372 = {_T_1371,wdata}; // @[Cat.scala 30:58:@3851.8]
  assign _GEN_69 = _T_604 ? {{1'd0}, _T_1372} : _GEN_68; // @[CSR.scala 278:29:@3849.6]
  assign _T_1374 = _T_336[31:0]; // @[CSR.scala 277:72:@3856.8]
  assign _T_1375 = {_T_1253,_T_1374}; // @[Cat.scala 30:58:@3857.8]
  assign _GEN_70 = _T_610 ? {{1'd0}, _T_1375} : _T_337; // @[CSR.scala 277:29:@3854.6]
  assign _T_1376 = _T_336[39:32]; // @[CSR.scala 278:45:@3861.8]
  assign _T_1377 = {_T_1376,wdata}; // @[Cat.scala 30:58:@3862.8]
  assign _GEN_71 = _T_608 ? {{1'd0}, _T_1377} : _GEN_70; // @[CSR.scala 278:29:@3860.6]
  assign _T_1379 = _T_339[31:0]; // @[CSR.scala 277:72:@3867.8]
  assign _T_1380 = {_T_1253,_T_1379}; // @[Cat.scala 30:58:@3868.8]
  assign _GEN_72 = _T_614 ? {{1'd0}, _T_1380} : _T_340; // @[CSR.scala 277:29:@3865.6]
  assign _T_1381 = _T_339[39:32]; // @[CSR.scala 278:45:@3872.8]
  assign _T_1382 = {_T_1381,wdata}; // @[Cat.scala 30:58:@3873.8]
  assign _GEN_73 = _T_612 ? {{1'd0}, _T_1382} : _GEN_72; // @[CSR.scala 278:29:@3871.6]
  assign _T_1384 = _T_342[31:0]; // @[CSR.scala 277:72:@3878.8]
  assign _T_1385 = {_T_1253,_T_1384}; // @[Cat.scala 30:58:@3879.8]
  assign _GEN_74 = _T_618 ? {{1'd0}, _T_1385} : _T_343; // @[CSR.scala 277:29:@3876.6]
  assign _T_1386 = _T_342[39:32]; // @[CSR.scala 278:45:@3883.8]
  assign _T_1387 = {_T_1386,wdata}; // @[Cat.scala 30:58:@3884.8]
  assign _GEN_75 = _T_616 ? {{1'd0}, _T_1387} : _GEN_74; // @[CSR.scala 278:29:@3882.6]
  assign _T_1389 = _T_345[31:0]; // @[CSR.scala 277:72:@3889.8]
  assign _T_1390 = {_T_1253,_T_1389}; // @[Cat.scala 30:58:@3890.8]
  assign _GEN_76 = _T_622 ? {{1'd0}, _T_1390} : _T_346; // @[CSR.scala 277:29:@3887.6]
  assign _T_1391 = _T_345[39:32]; // @[CSR.scala 278:45:@3894.8]
  assign _T_1392 = {_T_1391,wdata}; // @[Cat.scala 30:58:@3895.8]
  assign _GEN_77 = _T_620 ? {{1'd0}, _T_1392} : _GEN_76; // @[CSR.scala 278:29:@3893.6]
  assign _T_1394 = _T_348[31:0]; // @[CSR.scala 277:72:@3900.8]
  assign _T_1395 = {_T_1253,_T_1394}; // @[Cat.scala 30:58:@3901.8]
  assign _GEN_78 = _T_626 ? {{1'd0}, _T_1395} : _T_349; // @[CSR.scala 277:29:@3898.6]
  assign _T_1396 = _T_348[39:32]; // @[CSR.scala 278:45:@3905.8]
  assign _T_1397 = {_T_1396,wdata}; // @[Cat.scala 30:58:@3906.8]
  assign _GEN_79 = _T_624 ? {{1'd0}, _T_1397} : _GEN_78; // @[CSR.scala 278:29:@3904.6]
  assign _T_1399 = _T_351[31:0]; // @[CSR.scala 277:72:@3911.8]
  assign _T_1400 = {_T_1253,_T_1399}; // @[Cat.scala 30:58:@3912.8]
  assign _GEN_80 = _T_630 ? {{1'd0}, _T_1400} : _T_352; // @[CSR.scala 277:29:@3909.6]
  assign _T_1401 = _T_351[39:32]; // @[CSR.scala 278:45:@3916.8]
  assign _T_1402 = {_T_1401,wdata}; // @[Cat.scala 30:58:@3917.8]
  assign _GEN_81 = _T_628 ? {{1'd0}, _T_1402} : _GEN_80; // @[CSR.scala 278:29:@3915.6]
  assign _T_1404 = _T_354[31:0]; // @[CSR.scala 277:72:@3922.8]
  assign _T_1405 = {_T_1253,_T_1404}; // @[Cat.scala 30:58:@3923.8]
  assign _GEN_82 = _T_634 ? {{1'd0}, _T_1405} : _T_355; // @[CSR.scala 277:29:@3920.6]
  assign _T_1406 = _T_354[39:32]; // @[CSR.scala 278:45:@3927.8]
  assign _T_1407 = {_T_1406,wdata}; // @[Cat.scala 30:58:@3928.8]
  assign _GEN_83 = _T_632 ? {{1'd0}, _T_1407} : _GEN_82; // @[CSR.scala 278:29:@3926.6]
  assign _T_1409 = _T_357[31:0]; // @[CSR.scala 277:72:@3933.8]
  assign _T_1410 = {_T_1253,_T_1409}; // @[Cat.scala 30:58:@3934.8]
  assign _GEN_84 = _T_638 ? {{1'd0}, _T_1410} : _T_358; // @[CSR.scala 277:29:@3931.6]
  assign _T_1411 = _T_357[39:32]; // @[CSR.scala 278:45:@3938.8]
  assign _T_1412 = {_T_1411,wdata}; // @[Cat.scala 30:58:@3939.8]
  assign _GEN_85 = _T_636 ? {{1'd0}, _T_1412} : _GEN_84; // @[CSR.scala 278:29:@3937.6]
  assign _T_1414 = _T_249[31:0]; // @[CSR.scala 277:72:@3944.8]
  assign _T_1415 = {wdata,_T_1414}; // @[Cat.scala 30:58:@3945.8]
  assign _T_1416 = _T_1415[63:6]; // @[Util.scala 133:28:@3947.8]
  assign _GEN_86 = _T_640 ? _T_1415 : {{57'd0}, _T_241}; // @[CSR.scala 277:29:@3942.6]
  assign _GEN_87 = _T_640 ? _T_1416 : _GEN_0; // @[CSR.scala 277:29:@3942.6]
  assign _T_1417 = _T_249[63:32]; // @[CSR.scala 278:45:@3951.8]
  assign _T_1418 = {_T_1417,wdata}; // @[Cat.scala 30:58:@3952.8]
  assign _T_1419 = _T_1418[63:6]; // @[Util.scala 133:28:@3954.8]
  assign _GEN_88 = _T_478 ? _T_1418 : _GEN_86; // @[CSR.scala 278:29:@3950.6]
  assign _GEN_89 = _T_478 ? _T_1419 : _GEN_87; // @[CSR.scala 278:29:@3950.6]
  assign _T_1421 = _T_261[31:0]; // @[CSR.scala 277:72:@3959.8]
  assign _T_1422 = {wdata,_T_1421}; // @[Cat.scala 30:58:@3960.8]
  assign _T_1423 = _T_1422[63:6]; // @[Util.scala 133:28:@3962.8]
  assign _GEN_90 = _T_642 ? _T_1422 : {{57'd0}, _T_253}; // @[CSR.scala 277:29:@3957.6]
  assign _GEN_91 = _T_642 ? _T_1423 : _GEN_1; // @[CSR.scala 277:29:@3957.6]
  assign _T_1424 = _T_261[63:32]; // @[CSR.scala 278:45:@3966.8]
  assign _T_1425 = {_T_1424,wdata}; // @[Cat.scala 30:58:@3967.8]
  assign _T_1426 = _T_1425[63:6]; // @[Util.scala 133:28:@3969.8]
  assign _GEN_92 = _T_480 ? _T_1425 : _GEN_90; // @[CSR.scala 278:29:@3965.6]
  assign _GEN_93 = _T_480 ? _T_1426 : _GEN_91; // @[CSR.scala 278:29:@3965.6]
  assign _GEN_94 = _T_508 ? wdata : reg_dscratch; // @[CSR.scala 265:40:@3972.6]
  assign _T_1429 = wdata >> 2'h2; // @[CSR.scala 267:78:@3977.8]
  assign _GEN_225 = {{3'd0}, _T_1429}; // @[CSR.scala 267:86:@3978.8]
  assign _T_1431 = _GEN_225 << 2'h2; // @[CSR.scala 267:86:@3978.8]
  assign _GEN_95 = _T_500 ? _T_1431 : {{3'd0}, _GEN_15}; // @[CSR.scala 267:40:@3975.6]
  assign _GEN_96 = _T_498 ? wdata : reg_mscratch; // @[CSR.scala 268:40:@3981.6]
  assign _T_1433 = wdata & 32'h8000001f; // @[CSR.scala 269:62:@3985.8]
  assign _GEN_97 = _T_504 ? _T_1433 : _GEN_14; // @[CSR.scala 269:40:@3984.6]
  assign _GEN_98 = _T_502 ? wdata : _GEN_16; // @[CSR.scala 270:40:@3988.6]
  assign _GEN_99 = _T_510 ? wdata : reg_medeleg; // @[CSR.scala 271:42:@3992.6]
  assign _GEN_100 = wen ? _GEN_17 : _GEN_3; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_101 = wen ? _GEN_18 : _GEN_4; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_102 = wen ? _GEN_19 : reg_mip_msip; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_103 = wen ? _GEN_20 : reg_mie_msip; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_104 = wen ? _GEN_21 : reg_mie_mtip; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_105 = wen ? _GEN_23 : _T_265; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_106 = wen ? _GEN_25 : _T_268; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_107 = wen ? _GEN_27 : _T_271; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_108 = wen ? _GEN_29 : _T_274; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_109 = wen ? _GEN_31 : _T_277; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_110 = wen ? _GEN_33 : _T_280; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_111 = wen ? _GEN_35 : _T_283; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_112 = wen ? _GEN_37 : _T_286; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_113 = wen ? _GEN_39 : _T_289; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_114 = wen ? _GEN_41 : _T_292; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_115 = wen ? _GEN_43 : _T_295; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_116 = wen ? _GEN_45 : _T_298; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_117 = wen ? _GEN_47 : _T_301; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_118 = wen ? _GEN_49 : _T_304; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_119 = wen ? _GEN_51 : _T_307; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_120 = wen ? _GEN_53 : _T_310; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_121 = wen ? _GEN_55 : _T_313; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_122 = wen ? _GEN_57 : _T_316; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_123 = wen ? _GEN_59 : _T_319; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_124 = wen ? _GEN_61 : _T_322; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_125 = wen ? _GEN_63 : _T_325; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_126 = wen ? _GEN_65 : _T_328; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_127 = wen ? _GEN_67 : _T_331; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_128 = wen ? _GEN_69 : _T_334; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_129 = wen ? _GEN_71 : _T_337; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_130 = wen ? _GEN_73 : _T_340; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_131 = wen ? _GEN_75 : _T_343; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_132 = wen ? _GEN_77 : _T_346; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_133 = wen ? _GEN_79 : _T_349; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_134 = wen ? _GEN_81 : _T_352; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_135 = wen ? _GEN_83 : _T_355; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_136 = wen ? _GEN_85 : _T_358; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_137 = wen ? _GEN_88 : {{57'd0}, _T_241}; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_138 = wen ? _GEN_89 : _GEN_0; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_139 = wen ? _GEN_92 : {{57'd0}, _T_253}; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_140 = wen ? _GEN_93 : _GEN_1; // @[CSR.scala 242:14:@3521.4]
  assign _GEN_142 = wen ? _GEN_95 : {{3'd0}, _GEN_15}; // @[CSR.scala 242:14:@3521.4]
  assign io_rw_rdata = _T_1209[31:0]; // @[CSR.scala 240:15:@3520.4]
  assign io_eret = _T_940 | insn_ret; // @[CSR.scala 199:11:@3310.4]
  assign io_status_prv = reg_mstatus_prv; // @[CSR.scala 197:13:@3307.4]
  assign io_status_unimp5 = 14'h0; // @[CSR.scala 197:13:@3306.4]
  assign io_status_mprv = 1'h0; // @[CSR.scala 197:13:@3305.4]
  assign io_status_unimp4 = 2'h0; // @[CSR.scala 197:13:@3304.4]
  assign io_status_mpp = 2'h3; // @[CSR.scala 197:13:@3303.4]
  assign io_status_unimp3 = 3'h0; // @[CSR.scala 197:13:@3302.4]
  assign io_status_mpie = reg_mstatus_mpie; // @[CSR.scala 197:13:@3301.4]
  assign io_status_unimp2 = 3'h0; // @[CSR.scala 197:13:@3300.4]
  assign io_status_mie = reg_mstatus_mie; // @[CSR.scala 197:13:@3299.4]
  assign io_status_unimp1 = 3'h0; // @[CSR.scala 197:13:@3298.4]
  assign io_evec = io_xcpt ? 32'h80000004 : _GEN_10; // @[CSR.scala 212:13:@3331.6 CSR.scala 217:13:@3334.6 CSR.scala 224:13:@3341.6 CSR.scala 230:13:@3346.6]
  assign io_time = _T_249[31:0]; // @[CSR.scala 236:11:@3351.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_mstatus_prv = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  reg_mstatus_mpie = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  reg_mstatus_mie = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  reg_mepc = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  reg_mcause = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  reg_mtval = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  reg_mscratch = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  reg_medeleg = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  reg_mip_mtip = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  reg_mip_msip = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  reg_mie_mtip = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  reg_mie_msip = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_240 = _RAND_12[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {2{`RANDOM}};
  _T_244 = _RAND_13[57:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_252 = _RAND_14[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {2{`RANDOM}};
  _T_256 = _RAND_15[57:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {2{`RANDOM}};
  _T_264 = _RAND_16[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {2{`RANDOM}};
  _T_267 = _RAND_17[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {2{`RANDOM}};
  _T_270 = _RAND_18[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {2{`RANDOM}};
  _T_273 = _RAND_19[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {2{`RANDOM}};
  _T_276 = _RAND_20[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {2{`RANDOM}};
  _T_279 = _RAND_21[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {2{`RANDOM}};
  _T_282 = _RAND_22[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {2{`RANDOM}};
  _T_285 = _RAND_23[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {2{`RANDOM}};
  _T_288 = _RAND_24[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {2{`RANDOM}};
  _T_291 = _RAND_25[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {2{`RANDOM}};
  _T_294 = _RAND_26[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {2{`RANDOM}};
  _T_297 = _RAND_27[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {2{`RANDOM}};
  _T_300 = _RAND_28[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {2{`RANDOM}};
  _T_303 = _RAND_29[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {2{`RANDOM}};
  _T_306 = _RAND_30[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {2{`RANDOM}};
  _T_309 = _RAND_31[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {2{`RANDOM}};
  _T_312 = _RAND_32[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {2{`RANDOM}};
  _T_315 = _RAND_33[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {2{`RANDOM}};
  _T_318 = _RAND_34[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {2{`RANDOM}};
  _T_321 = _RAND_35[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {2{`RANDOM}};
  _T_324 = _RAND_36[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {2{`RANDOM}};
  _T_327 = _RAND_37[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {2{`RANDOM}};
  _T_330 = _RAND_38[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {2{`RANDOM}};
  _T_333 = _RAND_39[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {2{`RANDOM}};
  _T_336 = _RAND_40[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {2{`RANDOM}};
  _T_339 = _RAND_41[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {2{`RANDOM}};
  _T_342 = _RAND_42[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {2{`RANDOM}};
  _T_345 = _RAND_43[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {2{`RANDOM}};
  _T_348 = _RAND_44[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {2{`RANDOM}};
  _T_351 = _RAND_45[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {2{`RANDOM}};
  _T_354 = _RAND_46[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {2{`RANDOM}};
  _T_357 = _RAND_47[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  reg_dscratch = _RAND_48[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      reg_mstatus_prv <= 2'h3;
    end else begin
      if (_T_954) begin
        reg_mstatus_prv <= 2'h3;
      end
    end
    if (reset) begin
      reg_mstatus_mpie <= 1'h0;
    end else begin
      if (wen) begin
        if (_T_490) begin
          reg_mstatus_mpie <= _T_1222;
        end else begin
          if (_T_954) begin
            reg_mstatus_mpie <= 1'h1;
          end
        end
      end else begin
        if (_T_954) begin
          reg_mstatus_mpie <= 1'h1;
        end
      end
    end
    if (reset) begin
      reg_mstatus_mie <= 1'h0;
    end else begin
      if (wen) begin
        if (_T_490) begin
          reg_mstatus_mie <= _T_1220;
        end else begin
          if (_T_954) begin
            reg_mstatus_mie <= reg_mstatus_mpie;
          end
        end
      end else begin
        if (_T_954) begin
          reg_mstatus_mie <= reg_mstatus_mpie;
        end
      end
    end
    reg_mepc <= _GEN_142[31:0];
    if (wen) begin
      if (_T_504) begin
        reg_mcause <= _T_1433;
      end else begin
        if (io_xcpt) begin
          reg_mcause <= io_cause;
        end else begin
          if (insn_break) begin
            reg_mcause <= 32'h3;
          end else begin
            if (insn_call) begin
              reg_mcause <= {{28'd0}, _T_959};
            end
          end
        end
      end
    end else begin
      if (io_xcpt) begin
        reg_mcause <= io_cause;
      end else begin
        if (insn_break) begin
          reg_mcause <= 32'h3;
        end else begin
          if (insn_call) begin
            reg_mcause <= {{28'd0}, _T_959};
          end
        end
      end
    end
    if (wen) begin
      if (_T_502) begin
        reg_mtval <= wdata;
      end else begin
        if (io_xcpt) begin
          reg_mtval <= io_tval;
        end
      end
    end else begin
      if (io_xcpt) begin
        reg_mtval <= io_tval;
      end
    end
    if (wen) begin
      if (_T_498) begin
        reg_mscratch <= wdata;
      end
    end
    if (wen) begin
      if (_T_510) begin
        reg_medeleg <= wdata;
      end
    end
    if (reset) begin
      reg_mip_mtip <= 1'h0;
    end else begin
      reg_mip_mtip <= 1'h1;
    end
    if (reset) begin
      reg_mip_msip <= 1'h0;
    end else begin
      if (wen) begin
        if (_T_494) begin
          reg_mip_msip <= _T_1235;
        end
      end
    end
    if (reset) begin
      reg_mie_mtip <= 1'h0;
    end else begin
      if (wen) begin
        if (_T_496) begin
          reg_mie_mtip <= _T_1237;
        end
      end
    end
    if (reset) begin
      reg_mie_msip <= 1'h0;
    end else begin
      if (wen) begin
        if (_T_496) begin
          reg_mie_msip <= _T_1235;
        end
      end
    end
    if (reset) begin
      _T_240 <= 6'h0;
    end else begin
      _T_240 <= _GEN_137[5:0];
    end
    if (reset) begin
      _T_244 <= 58'h0;
    end else begin
      if (wen) begin
        if (_T_478) begin
          _T_244 <= _T_1419;
        end else begin
          if (_T_640) begin
            _T_244 <= _T_1416;
          end else begin
            if (_T_245) begin
              _T_244 <= _T_248;
            end
          end
        end
      end else begin
        if (_T_245) begin
          _T_244 <= _T_248;
        end
      end
    end
    if (reset) begin
      _T_252 <= 6'h0;
    end else begin
      _T_252 <= _GEN_139[5:0];
    end
    if (reset) begin
      _T_256 <= 58'h0;
    end else begin
      if (wen) begin
        if (_T_480) begin
          _T_256 <= _T_1426;
        end else begin
          if (_T_642) begin
            _T_256 <= _T_1423;
          end else begin
            if (_T_257) begin
              _T_256 <= _T_260;
            end
          end
        end
      end else begin
        if (_T_257) begin
          _T_256 <= _T_260;
        end
      end
    end
    _T_264 <= _GEN_105[39:0];
    _T_267 <= _GEN_106[39:0];
    _T_270 <= _GEN_107[39:0];
    _T_273 <= _GEN_108[39:0];
    _T_276 <= _GEN_109[39:0];
    _T_279 <= _GEN_110[39:0];
    _T_282 <= _GEN_111[39:0];
    _T_285 <= _GEN_112[39:0];
    _T_288 <= _GEN_113[39:0];
    _T_291 <= _GEN_114[39:0];
    _T_294 <= _GEN_115[39:0];
    _T_297 <= _GEN_116[39:0];
    _T_300 <= _GEN_117[39:0];
    _T_303 <= _GEN_118[39:0];
    _T_306 <= _GEN_119[39:0];
    _T_309 <= _GEN_120[39:0];
    _T_312 <= _GEN_121[39:0];
    _T_315 <= _GEN_122[39:0];
    _T_318 <= _GEN_123[39:0];
    _T_321 <= _GEN_124[39:0];
    _T_324 <= _GEN_125[39:0];
    _T_327 <= _GEN_126[39:0];
    _T_330 <= _GEN_127[39:0];
    _T_333 <= _GEN_128[39:0];
    _T_336 <= _GEN_129[39:0];
    _T_339 <= _GEN_130[39:0];
    _T_342 <= _GEN_131[39:0];
    _T_345 <= _GEN_132[39:0];
    _T_348 <= _GEN_133[39:0];
    _T_351 <= _GEN_134[39:0];
    _T_354 <= _GEN_135[39:0];
    _T_357 <= _GEN_136[39:0];
    if (wen) begin
      if (_T_508) begin
        reg_dscratch <= wdata;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_948) begin
          $fwrite(32'h80000002,"Assertion failed: these conditions must be mutually exclusive\n    at CSR.scala:201 assert(PopCount(insn_ret :: io.illegal :: Nil) <= 1, \"these conditions must be mutually exclusive\")\n"); // @[CSR.scala 201:9:@3317.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_948) begin
          $fatal; // @[CSR.scala 201:9:@3318.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
