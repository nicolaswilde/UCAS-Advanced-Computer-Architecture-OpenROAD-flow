module ALU( // @[:@4914.2]
  input  [31:0] io_op1, // @[:@4917.4]
  input  [31:0] io_op2, // @[:@4917.4]
  input  [31:0] io_pc, // @[:@4917.4]
  input  [3:0]  io_ctrl_fun, // @[:@4917.4]
  input  [3:0]  io_ctrl_br_type, // @[:@4917.4]
  input  [1:0]  io_ctrl_wb_sel, // @[:@4917.4]
  output [1:0]  io_ctrl_pc_sel, // @[:@4917.4]
  input  [31:0] io_rs2_data, // @[:@4917.4]
  output [31:0] io_result, // @[:@4917.4]
  output [31:0] io_target_brjmp, // @[:@4917.4]
  output [31:0] io_target_jpreg, // @[:@4917.4]
  output [31:0] io_target_conti // @[:@4917.4]
);
  wire [4:0] alu_shamt; // @[ALU.scala 32:32:@4919.4]
  wire [32:0] _T_25; // @[ALU.scala 33:34:@4920.4]
  wire [31:0] add_result; // @[ALU.scala 33:34:@4921.4]
  wire  _T_29; // @[ALU.scala 38:18:@4924.4]
  wire  _T_30; // @[ALU.scala 39:18:@4925.4]
  wire [32:0] _T_31; // @[ALU.scala 39:44:@4926.4]
  wire [32:0] _T_32; // @[ALU.scala 39:44:@4927.4]
  wire [31:0] _T_33; // @[ALU.scala 39:44:@4928.4]
  wire  _T_34; // @[ALU.scala 40:18:@4929.4]
  wire [31:0] _T_35; // @[ALU.scala 40:44:@4930.4]
  wire  _T_36; // @[ALU.scala 41:18:@4931.4]
  wire [31:0] _T_37; // @[ALU.scala 41:44:@4932.4]
  wire  _T_38; // @[ALU.scala 42:18:@4933.4]
  wire [31:0] _T_39; // @[ALU.scala 42:44:@4934.4]
  wire  _T_40; // @[ALU.scala 43:18:@4935.4]
  wire [31:0] _T_41; // @[ALU.scala 43:44:@4936.4]
  wire [31:0] _T_42; // @[ALU.scala 43:60:@4937.4]
  wire  _T_43; // @[ALU.scala 43:51:@4938.4]
  wire  _T_44; // @[ALU.scala 44:18:@4939.4]
  wire  _T_45; // @[ALU.scala 44:44:@4940.4]
  wire  _T_46; // @[ALU.scala 45:18:@4941.4]
  wire [62:0] _GEN_0; // @[ALU.scala 45:44:@4942.4]
  wire [62:0] _T_47; // @[ALU.scala 45:44:@4942.4]
  wire [31:0] _T_48; // @[ALU.scala 45:57:@4943.4]
  wire  _T_49; // @[ALU.scala 46:18:@4944.4]
  wire [31:0] _T_51; // @[ALU.scala 46:51:@4946.4]
  wire [31:0] _T_52; // @[ALU.scala 46:65:@4947.4]
  wire  _T_53; // @[ALU.scala 47:18:@4948.4]
  wire [31:0] _T_54; // @[ALU.scala 47:44:@4949.4]
  wire  _T_55; // @[ALU.scala 48:18:@4950.4]
  wire  _T_56; // @[ALU.scala 49:18:@4951.4]
  wire [31:0] _T_57; // @[Mux.scala 61:16:@4952.4]
  wire [31:0] _T_58; // @[Mux.scala 61:16:@4953.4]
  wire [31:0] _T_59; // @[Mux.scala 61:16:@4954.4]
  wire [31:0] _T_60; // @[Mux.scala 61:16:@4955.4]
  wire [31:0] _T_61; // @[Mux.scala 61:16:@4956.4]
  wire [31:0] _T_62; // @[Mux.scala 61:16:@4957.4]
  wire [31:0] _T_63; // @[Mux.scala 61:16:@4958.4]
  wire [31:0] _T_64; // @[Mux.scala 61:16:@4959.4]
  wire [31:0] _T_65; // @[Mux.scala 61:16:@4960.4]
  wire [31:0] _T_66; // @[Mux.scala 61:16:@4961.4]
  wire [31:0] _T_67; // @[Mux.scala 61:16:@4962.4]
  wire [31:0] result; // @[Mux.scala 61:16:@4963.4]
  wire [32:0] _T_69; // @[ALU.scala 52:31:@4965.4]
  wire [30:0] _T_71; // @[ALU.scala 53:39:@4968.4]
  wire [32:0] _T_75; // @[ALU.scala 54:31:@4971.4]
  wire  _T_77; // @[ALU.scala 55:40:@4974.4]
  wire  br_eq; // @[ALU.scala 57:29:@4977.4]
  wire [31:0] _T_80; // @[ALU.scala 58:50:@4979.4]
  wire  br_lt; // @[ALU.scala 58:36:@4980.4]
  wire  br_ltu; // @[ALU.scala 59:36:@4981.4]
  wire  _T_81; // @[ALU.scala 63:25:@4982.4]
  wire  _T_82; // @[ALU.scala 64:25:@4983.4]
  wire  _T_84; // @[ALU.scala 64:41:@4984.4]
  wire [1:0] _T_85; // @[ALU.scala 64:40:@4985.4]
  wire  _T_86; // @[ALU.scala 65:25:@4986.4]
  wire [1:0] _T_87; // @[ALU.scala 65:40:@4987.4]
  wire  _T_88; // @[ALU.scala 66:25:@4988.4]
  wire  _T_90; // @[ALU.scala 66:41:@4989.4]
  wire [1:0] _T_91; // @[ALU.scala 66:40:@4990.4]
  wire  _T_92; // @[ALU.scala 67:25:@4991.4]
  wire  _T_94; // @[ALU.scala 67:41:@4992.4]
  wire [1:0] _T_95; // @[ALU.scala 67:40:@4993.4]
  wire  _T_96; // @[ALU.scala 68:25:@4994.4]
  wire [1:0] _T_97; // @[ALU.scala 68:40:@4995.4]
  wire  _T_98; // @[ALU.scala 69:25:@4996.4]
  wire [1:0] _T_99; // @[ALU.scala 69:40:@4997.4]
  wire  _T_100; // @[ALU.scala 70:25:@4998.4]
  wire  _T_101; // @[ALU.scala 71:25:@4999.4]
  wire [1:0] _T_102; // @[ALU.scala 71:8:@5000.4]
  wire [1:0] _T_103; // @[ALU.scala 70:8:@5001.4]
  wire [1:0] _T_104; // @[ALU.scala 69:8:@5002.4]
  wire [1:0] _T_105; // @[ALU.scala 68:8:@5003.4]
  wire [1:0] _T_106; // @[ALU.scala 67:8:@5004.4]
  wire [1:0] _T_107; // @[ALU.scala 66:8:@5005.4]
  wire [1:0] _T_108; // @[ALU.scala 65:8:@5006.4]
  wire [1:0] _T_109; // @[ALU.scala 64:8:@5007.4]
  assign alu_shamt = io_op2[4:0]; // @[ALU.scala 32:32:@4919.4]
  assign _T_25 = io_op1 + io_op2; // @[ALU.scala 33:34:@4920.4]
  assign add_result = io_op1 + io_op2; // @[ALU.scala 33:34:@4921.4]
  assign _T_29 = io_ctrl_fun == 4'h0; // @[ALU.scala 38:18:@4924.4]
  assign _T_30 = io_ctrl_fun == 4'h1; // @[ALU.scala 39:18:@4925.4]
  assign _T_31 = io_op1 - io_op2; // @[ALU.scala 39:44:@4926.4]
  assign _T_32 = $unsigned(_T_31); // @[ALU.scala 39:44:@4927.4]
  assign _T_33 = _T_32[31:0]; // @[ALU.scala 39:44:@4928.4]
  assign _T_34 = io_ctrl_fun == 4'h5; // @[ALU.scala 40:18:@4929.4]
  assign _T_35 = io_op1 & io_op2; // @[ALU.scala 40:44:@4930.4]
  assign _T_36 = io_ctrl_fun == 4'h6; // @[ALU.scala 41:18:@4931.4]
  assign _T_37 = io_op1 | io_op2; // @[ALU.scala 41:44:@4932.4]
  assign _T_38 = io_ctrl_fun == 4'h7; // @[ALU.scala 42:18:@4933.4]
  assign _T_39 = io_op1 ^ io_op2; // @[ALU.scala 42:44:@4934.4]
  assign _T_40 = io_ctrl_fun == 4'h8; // @[ALU.scala 43:18:@4935.4]
  assign _T_41 = $signed(io_op1); // @[ALU.scala 43:44:@4936.4]
  assign _T_42 = $signed(io_op2); // @[ALU.scala 43:60:@4937.4]
  assign _T_43 = $signed(_T_41) < $signed(_T_42); // @[ALU.scala 43:51:@4938.4]
  assign _T_44 = io_ctrl_fun == 4'h9; // @[ALU.scala 44:18:@4939.4]
  assign _T_45 = io_op1 < io_op2; // @[ALU.scala 44:44:@4940.4]
  assign _T_46 = io_ctrl_fun == 4'h2; // @[ALU.scala 45:18:@4941.4]
  assign _GEN_0 = {{31'd0}, io_op1}; // @[ALU.scala 45:44:@4942.4]
  assign _T_47 = _GEN_0 << alu_shamt; // @[ALU.scala 45:44:@4942.4]
  assign _T_48 = _T_47[31:0]; // @[ALU.scala 45:57:@4943.4]
  assign _T_49 = io_ctrl_fun == 4'h4; // @[ALU.scala 46:18:@4944.4]
  assign _T_51 = $signed(_T_41) >>> alu_shamt; // @[ALU.scala 46:51:@4946.4]
  assign _T_52 = $unsigned(_T_51); // @[ALU.scala 46:65:@4947.4]
  assign _T_53 = io_ctrl_fun == 4'h3; // @[ALU.scala 47:18:@4948.4]
  assign _T_54 = io_op1 >> alu_shamt; // @[ALU.scala 47:44:@4949.4]
  assign _T_55 = io_ctrl_fun == 4'ha; // @[ALU.scala 48:18:@4950.4]
  assign _T_56 = io_ctrl_fun == 4'hb; // @[ALU.scala 49:18:@4951.4]
  assign _T_57 = _T_56 ? io_op2 : 32'h0; // @[Mux.scala 61:16:@4952.4]
  assign _T_58 = _T_55 ? io_op1 : _T_57; // @[Mux.scala 61:16:@4953.4]
  assign _T_59 = _T_53 ? _T_54 : _T_58; // @[Mux.scala 61:16:@4954.4]
  assign _T_60 = _T_49 ? _T_52 : _T_59; // @[Mux.scala 61:16:@4955.4]
  assign _T_61 = _T_46 ? _T_48 : _T_60; // @[Mux.scala 61:16:@4956.4]
  assign _T_62 = _T_44 ? {{31'd0}, _T_45} : _T_61; // @[Mux.scala 61:16:@4957.4]
  assign _T_63 = _T_40 ? {{31'd0}, _T_43} : _T_62; // @[Mux.scala 61:16:@4958.4]
  assign _T_64 = _T_38 ? _T_39 : _T_63; // @[Mux.scala 61:16:@4959.4]
  assign _T_65 = _T_36 ? _T_37 : _T_64; // @[Mux.scala 61:16:@4960.4]
  assign _T_66 = _T_34 ? _T_35 : _T_65; // @[Mux.scala 61:16:@4961.4]
  assign _T_67 = _T_30 ? _T_33 : _T_66; // @[Mux.scala 61:16:@4962.4]
  assign result = _T_29 ? add_result : _T_67; // @[Mux.scala 61:16:@4963.4]
  assign _T_69 = io_pc + io_op2; // @[ALU.scala 52:31:@4965.4]
  assign _T_71 = add_result[31:1]; // @[ALU.scala 53:39:@4968.4]
  assign _T_75 = io_pc + 32'h4; // @[ALU.scala 54:31:@4971.4]
  assign _T_77 = io_ctrl_wb_sel == 2'h2; // @[ALU.scala 55:40:@4974.4]
  assign br_eq = io_op1 == io_rs2_data; // @[ALU.scala 57:29:@4977.4]
  assign _T_80 = $signed(io_rs2_data); // @[ALU.scala 58:50:@4979.4]
  assign br_lt = $signed(_T_41) < $signed(_T_80); // @[ALU.scala 58:36:@4980.4]
  assign br_ltu = io_op1 < io_rs2_data; // @[ALU.scala 59:36:@4981.4]
  assign _T_81 = io_ctrl_br_type == 4'h0; // @[ALU.scala 63:25:@4982.4]
  assign _T_82 = io_ctrl_br_type == 4'h1; // @[ALU.scala 64:25:@4983.4]
  assign _T_84 = br_eq == 1'h0; // @[ALU.scala 64:41:@4984.4]
  assign _T_85 = _T_84 ? 2'h1 : 2'h0; // @[ALU.scala 64:40:@4985.4]
  assign _T_86 = io_ctrl_br_type == 4'h2; // @[ALU.scala 65:25:@4986.4]
  assign _T_87 = br_eq ? 2'h1 : 2'h0; // @[ALU.scala 65:40:@4987.4]
  assign _T_88 = io_ctrl_br_type == 4'h3; // @[ALU.scala 66:25:@4988.4]
  assign _T_90 = br_lt == 1'h0; // @[ALU.scala 66:41:@4989.4]
  assign _T_91 = _T_90 ? 2'h1 : 2'h0; // @[ALU.scala 66:40:@4990.4]
  assign _T_92 = io_ctrl_br_type == 4'h4; // @[ALU.scala 67:25:@4991.4]
  assign _T_94 = br_ltu == 1'h0; // @[ALU.scala 67:41:@4992.4]
  assign _T_95 = _T_94 ? 2'h1 : 2'h0; // @[ALU.scala 67:40:@4993.4]
  assign _T_96 = io_ctrl_br_type == 4'h5; // @[ALU.scala 68:25:@4994.4]
  assign _T_97 = br_lt ? 2'h1 : 2'h0; // @[ALU.scala 68:40:@4995.4]
  assign _T_98 = io_ctrl_br_type == 4'h6; // @[ALU.scala 69:25:@4996.4]
  assign _T_99 = br_ltu ? 2'h1 : 2'h0; // @[ALU.scala 69:40:@4997.4]
  assign _T_100 = io_ctrl_br_type == 4'h7; // @[ALU.scala 70:25:@4998.4]
  assign _T_101 = io_ctrl_br_type == 4'h8; // @[ALU.scala 71:25:@4999.4]
  assign _T_102 = _T_101 ? 2'h2 : 2'h0; // @[ALU.scala 71:8:@5000.4]
  assign _T_103 = _T_100 ? 2'h1 : _T_102; // @[ALU.scala 70:8:@5001.4]
  assign _T_104 = _T_98 ? _T_99 : _T_103; // @[ALU.scala 69:8:@5002.4]
  assign _T_105 = _T_96 ? _T_97 : _T_104; // @[ALU.scala 68:8:@5003.4]
  assign _T_106 = _T_92 ? _T_95 : _T_105; // @[ALU.scala 67:8:@5004.4]
  assign _T_107 = _T_88 ? _T_91 : _T_106; // @[ALU.scala 66:8:@5005.4]
  assign _T_108 = _T_86 ? _T_87 : _T_107; // @[ALU.scala 65:8:@5006.4]
  assign _T_109 = _T_82 ? _T_85 : _T_108; // @[ALU.scala 64:8:@5007.4]
  assign io_ctrl_pc_sel = _T_81 ? 2'h0 : _T_109; // @[ALU.scala 62:18:@5009.4]
  assign io_result = _T_77 ? io_target_conti : result; // @[ALU.scala 55:18:@4976.4]
  assign io_target_brjmp = io_pc + io_op2; // @[ALU.scala 52:22:@4967.4]
  assign io_target_jpreg = {_T_71,1'h0}; // @[ALU.scala 53:22:@4970.4]
  assign io_target_conti = io_pc + 32'h4; // @[ALU.scala 54:22:@4973.4]
endmodule
