module InstDecoder( // @[:@3996.2]
  input  [31:0] io_inst, // @[:@3999.4]
  output [3:0]  io_cinfo_br_type, // @[:@3999.4]
  output [1:0]  io_cinfo_op1_sel, // @[:@3999.4]
  output [2:0]  io_cinfo_op2_sel, // @[:@3999.4]
  output        io_cinfo_rs1_oen, // @[:@3999.4]
  output        io_cinfo_rs2_oen, // @[:@3999.4]
  output [3:0]  io_cinfo_alu_fun, // @[:@3999.4]
  output [1:0]  io_cinfo_wb_sel, // @[:@3999.4]
  output        io_cinfo_rf_wen, // @[:@3999.4]
  output        io_cinfo_mem_en, // @[:@3999.4]
  output        io_cinfo_mem_fcn, // @[:@3999.4]
  output [2:0]  io_cinfo_mem_typ, // @[:@3999.4]
  output [2:0]  io_cinfo_csr_cmd, // @[:@3999.4]
  output        io_cinfo_illegal, // @[:@3999.4]
  output        io_cinfo_fencei, // @[:@3999.4]
  output        io_cinfo_is_branch, // @[:@3999.4]
  output        io_cinfo_push, // @[:@3999.4]
  output        io_cinfo_pop, // @[:@3999.4]
  output [4:0]  io_cinfo_rs1_addr, // @[:@3999.4]
  output [4:0]  io_cinfo_rs2_addr, // @[:@3999.4]
  output [4:0]  io_cinfo_wbaddr, // @[:@3999.4]
  output [31:0] io_dinfo_imm_i, // @[:@3999.4]
  output [31:0] io_dinfo_imm_s, // @[:@3999.4]
  output [31:0] io_dinfo_imm_sb, // @[:@3999.4]
  output [31:0] io_dinfo_imm_u, // @[:@3999.4]
  output [31:0] io_dinfo_imm_uj, // @[:@3999.4]
  output [31:0] io_dinfo_imm_z // @[:@3999.4]
);
  wire [31:0] _T_13; // @[Lookup.scala 9:38:@4001.4]
  wire  _T_14; // @[Lookup.scala 9:38:@4002.4]
  wire  _T_18; // @[Lookup.scala 9:38:@4004.4]
  wire  _T_22; // @[Lookup.scala 9:38:@4006.4]
  wire  _T_26; // @[Lookup.scala 9:38:@4008.4]
  wire  _T_30; // @[Lookup.scala 9:38:@4010.4]
  wire  _T_34; // @[Lookup.scala 9:38:@4012.4]
  wire  _T_38; // @[Lookup.scala 9:38:@4014.4]
  wire  _T_42; // @[Lookup.scala 9:38:@4016.4]
  wire [31:0] _T_45; // @[Lookup.scala 9:38:@4017.4]
  wire  _T_46; // @[Lookup.scala 9:38:@4018.4]
  wire  _T_50; // @[Lookup.scala 9:38:@4020.4]
  wire  _T_54; // @[Lookup.scala 9:38:@4022.4]
  wire  _T_58; // @[Lookup.scala 9:38:@4024.4]
  wire  _T_62; // @[Lookup.scala 9:38:@4026.4]
  wire  _T_66; // @[Lookup.scala 9:38:@4028.4]
  wire  _T_70; // @[Lookup.scala 9:38:@4030.4]
  wire  _T_74; // @[Lookup.scala 9:38:@4032.4]
  wire [31:0] _T_77; // @[Lookup.scala 9:38:@4033.4]
  wire  _T_78; // @[Lookup.scala 9:38:@4034.4]
  wire  _T_82; // @[Lookup.scala 9:38:@4036.4]
  wire  _T_86; // @[Lookup.scala 9:38:@4038.4]
  wire [31:0] _T_89; // @[Lookup.scala 9:38:@4039.4]
  wire  _T_90; // @[Lookup.scala 9:38:@4040.4]
  wire  _T_94; // @[Lookup.scala 9:38:@4042.4]
  wire  _T_98; // @[Lookup.scala 9:38:@4044.4]
  wire  _T_102; // @[Lookup.scala 9:38:@4046.4]
  wire  _T_106; // @[Lookup.scala 9:38:@4048.4]
  wire  _T_110; // @[Lookup.scala 9:38:@4050.4]
  wire  _T_114; // @[Lookup.scala 9:38:@4052.4]
  wire  _T_118; // @[Lookup.scala 9:38:@4054.4]
  wire  _T_122; // @[Lookup.scala 9:38:@4056.4]
  wire  _T_126; // @[Lookup.scala 9:38:@4058.4]
  wire  _T_130; // @[Lookup.scala 9:38:@4060.4]
  wire  _T_134; // @[Lookup.scala 9:38:@4062.4]
  wire  _T_138; // @[Lookup.scala 9:38:@4064.4]
  wire  _T_142; // @[Lookup.scala 9:38:@4066.4]
  wire  _T_146; // @[Lookup.scala 9:38:@4068.4]
  wire  _T_150; // @[Lookup.scala 9:38:@4070.4]
  wire  _T_154; // @[Lookup.scala 9:38:@4072.4]
  wire  _T_158; // @[Lookup.scala 9:38:@4074.4]
  wire  _T_162; // @[Lookup.scala 9:38:@4076.4]
  wire  _T_166; // @[Lookup.scala 9:38:@4078.4]
  wire  _T_170; // @[Lookup.scala 9:38:@4080.4]
  wire  _T_174; // @[Lookup.scala 9:38:@4082.4]
  wire  _T_178; // @[Lookup.scala 9:38:@4084.4]
  wire  _T_182; // @[Lookup.scala 9:38:@4086.4]
  wire  _T_186; // @[Lookup.scala 9:38:@4088.4]
  wire  _T_190; // @[Lookup.scala 9:38:@4090.4]
  wire  _T_194; // @[Lookup.scala 9:38:@4092.4]
  wire  _T_198; // @[Lookup.scala 9:38:@4094.4]
  wire  _T_202; // @[Lookup.scala 9:38:@4096.4]
  wire  _T_206; // @[Lookup.scala 9:38:@4098.4]
  wire  _T_210; // @[Lookup.scala 9:38:@4100.4]
  wire  _T_212; // @[Lookup.scala 11:37:@4102.4]
  wire  _T_213; // @[Lookup.scala 11:37:@4103.4]
  wire  _T_214; // @[Lookup.scala 11:37:@4104.4]
  wire  _T_215; // @[Lookup.scala 11:37:@4105.4]
  wire  _T_216; // @[Lookup.scala 11:37:@4106.4]
  wire  _T_217; // @[Lookup.scala 11:37:@4107.4]
  wire  _T_218; // @[Lookup.scala 11:37:@4108.4]
  wire  _T_219; // @[Lookup.scala 11:37:@4109.4]
  wire  _T_220; // @[Lookup.scala 11:37:@4110.4]
  wire  _T_221; // @[Lookup.scala 11:37:@4111.4]
  wire  _T_222; // @[Lookup.scala 11:37:@4112.4]
  wire  _T_223; // @[Lookup.scala 11:37:@4113.4]
  wire  _T_224; // @[Lookup.scala 11:37:@4114.4]
  wire  _T_225; // @[Lookup.scala 11:37:@4115.4]
  wire  _T_226; // @[Lookup.scala 11:37:@4116.4]
  wire  _T_227; // @[Lookup.scala 11:37:@4117.4]
  wire  _T_228; // @[Lookup.scala 11:37:@4118.4]
  wire  _T_229; // @[Lookup.scala 11:37:@4119.4]
  wire  _T_230; // @[Lookup.scala 11:37:@4120.4]
  wire  _T_231; // @[Lookup.scala 11:37:@4121.4]
  wire  _T_232; // @[Lookup.scala 11:37:@4122.4]
  wire  _T_233; // @[Lookup.scala 11:37:@4123.4]
  wire  _T_234; // @[Lookup.scala 11:37:@4124.4]
  wire  _T_235; // @[Lookup.scala 11:37:@4125.4]
  wire  _T_236; // @[Lookup.scala 11:37:@4126.4]
  wire  _T_237; // @[Lookup.scala 11:37:@4127.4]
  wire  _T_238; // @[Lookup.scala 11:37:@4128.4]
  wire  _T_239; // @[Lookup.scala 11:37:@4129.4]
  wire  _T_240; // @[Lookup.scala 11:37:@4130.4]
  wire  _T_241; // @[Lookup.scala 11:37:@4131.4]
  wire  _T_242; // @[Lookup.scala 11:37:@4132.4]
  wire  _T_243; // @[Lookup.scala 11:37:@4133.4]
  wire  _T_244; // @[Lookup.scala 11:37:@4134.4]
  wire  _T_245; // @[Lookup.scala 11:37:@4135.4]
  wire  _T_246; // @[Lookup.scala 11:37:@4136.4]
  wire  _T_247; // @[Lookup.scala 11:37:@4137.4]
  wire  _T_248; // @[Lookup.scala 11:37:@4138.4]
  wire  _T_249; // @[Lookup.scala 11:37:@4139.4]
  wire  _T_250; // @[Lookup.scala 11:37:@4140.4]
  wire  _T_251; // @[Lookup.scala 11:37:@4141.4]
  wire  _T_252; // @[Lookup.scala 11:37:@4142.4]
  wire  _T_253; // @[Lookup.scala 11:37:@4143.4]
  wire  _T_254; // @[Lookup.scala 11:37:@4144.4]
  wire  _T_255; // @[Lookup.scala 11:37:@4145.4]
  wire  _T_256; // @[Lookup.scala 11:37:@4146.4]
  wire  _T_257; // @[Lookup.scala 11:37:@4147.4]
  wire  _T_258; // @[Lookup.scala 11:37:@4148.4]
  wire  _T_259; // @[Lookup.scala 11:37:@4149.4]
  wire  signals_0; // @[Lookup.scala 11:37:@4150.4]
  wire [3:0] _T_273; // @[Lookup.scala 11:37:@4164.4]
  wire [3:0] _T_274; // @[Lookup.scala 11:37:@4165.4]
  wire [3:0] _T_275; // @[Lookup.scala 11:37:@4166.4]
  wire [3:0] _T_276; // @[Lookup.scala 11:37:@4167.4]
  wire [3:0] _T_277; // @[Lookup.scala 11:37:@4168.4]
  wire [3:0] _T_278; // @[Lookup.scala 11:37:@4169.4]
  wire [3:0] _T_279; // @[Lookup.scala 11:37:@4170.4]
  wire [3:0] _T_280; // @[Lookup.scala 11:37:@4171.4]
  wire [3:0] _T_281; // @[Lookup.scala 11:37:@4172.4]
  wire [3:0] _T_282; // @[Lookup.scala 11:37:@4173.4]
  wire [3:0] _T_283; // @[Lookup.scala 11:37:@4174.4]
  wire [3:0] _T_284; // @[Lookup.scala 11:37:@4175.4]
  wire [3:0] _T_285; // @[Lookup.scala 11:37:@4176.4]
  wire [3:0] _T_286; // @[Lookup.scala 11:37:@4177.4]
  wire [3:0] _T_287; // @[Lookup.scala 11:37:@4178.4]
  wire [3:0] _T_288; // @[Lookup.scala 11:37:@4179.4]
  wire [3:0] _T_289; // @[Lookup.scala 11:37:@4180.4]
  wire [3:0] _T_290; // @[Lookup.scala 11:37:@4181.4]
  wire [3:0] _T_291; // @[Lookup.scala 11:37:@4182.4]
  wire [3:0] _T_292; // @[Lookup.scala 11:37:@4183.4]
  wire [3:0] _T_293; // @[Lookup.scala 11:37:@4184.4]
  wire [3:0] _T_294; // @[Lookup.scala 11:37:@4185.4]
  wire [3:0] _T_295; // @[Lookup.scala 11:37:@4186.4]
  wire [3:0] _T_296; // @[Lookup.scala 11:37:@4187.4]
  wire [3:0] _T_297; // @[Lookup.scala 11:37:@4188.4]
  wire [3:0] _T_298; // @[Lookup.scala 11:37:@4189.4]
  wire [3:0] _T_299; // @[Lookup.scala 11:37:@4190.4]
  wire [3:0] _T_300; // @[Lookup.scala 11:37:@4191.4]
  wire [3:0] _T_301; // @[Lookup.scala 11:37:@4192.4]
  wire [3:0] _T_302; // @[Lookup.scala 11:37:@4193.4]
  wire [3:0] _T_303; // @[Lookup.scala 11:37:@4194.4]
  wire [3:0] _T_304; // @[Lookup.scala 11:37:@4195.4]
  wire [3:0] _T_305; // @[Lookup.scala 11:37:@4196.4]
  wire [3:0] _T_306; // @[Lookup.scala 11:37:@4197.4]
  wire [3:0] _T_307; // @[Lookup.scala 11:37:@4198.4]
  wire [3:0] _T_308; // @[Lookup.scala 11:37:@4199.4]
  wire [1:0] _T_316; // @[Lookup.scala 11:37:@4208.4]
  wire [1:0] _T_317; // @[Lookup.scala 11:37:@4209.4]
  wire [1:0] _T_318; // @[Lookup.scala 11:37:@4210.4]
  wire [1:0] _T_319; // @[Lookup.scala 11:37:@4211.4]
  wire [1:0] _T_320; // @[Lookup.scala 11:37:@4212.4]
  wire [1:0] _T_321; // @[Lookup.scala 11:37:@4213.4]
  wire [1:0] _T_322; // @[Lookup.scala 11:37:@4214.4]
  wire [1:0] _T_323; // @[Lookup.scala 11:37:@4215.4]
  wire [1:0] _T_324; // @[Lookup.scala 11:37:@4216.4]
  wire [1:0] _T_325; // @[Lookup.scala 11:37:@4217.4]
  wire [1:0] _T_326; // @[Lookup.scala 11:37:@4218.4]
  wire [1:0] _T_327; // @[Lookup.scala 11:37:@4219.4]
  wire [1:0] _T_328; // @[Lookup.scala 11:37:@4220.4]
  wire [1:0] _T_329; // @[Lookup.scala 11:37:@4221.4]
  wire [1:0] _T_330; // @[Lookup.scala 11:37:@4222.4]
  wire [1:0] _T_331; // @[Lookup.scala 11:37:@4223.4]
  wire [1:0] _T_332; // @[Lookup.scala 11:37:@4224.4]
  wire [1:0] _T_333; // @[Lookup.scala 11:37:@4225.4]
  wire [1:0] _T_334; // @[Lookup.scala 11:37:@4226.4]
  wire [1:0] _T_335; // @[Lookup.scala 11:37:@4227.4]
  wire [1:0] _T_336; // @[Lookup.scala 11:37:@4228.4]
  wire [1:0] _T_337; // @[Lookup.scala 11:37:@4229.4]
  wire [1:0] _T_338; // @[Lookup.scala 11:37:@4230.4]
  wire [1:0] _T_339; // @[Lookup.scala 11:37:@4231.4]
  wire [1:0] _T_340; // @[Lookup.scala 11:37:@4232.4]
  wire [1:0] _T_341; // @[Lookup.scala 11:37:@4233.4]
  wire [1:0] _T_342; // @[Lookup.scala 11:37:@4234.4]
  wire [1:0] _T_343; // @[Lookup.scala 11:37:@4235.4]
  wire [1:0] _T_344; // @[Lookup.scala 11:37:@4236.4]
  wire [1:0] _T_345; // @[Lookup.scala 11:37:@4237.4]
  wire [1:0] _T_346; // @[Lookup.scala 11:37:@4238.4]
  wire [1:0] _T_347; // @[Lookup.scala 11:37:@4239.4]
  wire [1:0] _T_348; // @[Lookup.scala 11:37:@4240.4]
  wire [1:0] _T_349; // @[Lookup.scala 11:37:@4241.4]
  wire [1:0] _T_350; // @[Lookup.scala 11:37:@4242.4]
  wire [1:0] _T_351; // @[Lookup.scala 11:37:@4243.4]
  wire [1:0] _T_352; // @[Lookup.scala 11:37:@4244.4]
  wire [1:0] _T_353; // @[Lookup.scala 11:37:@4245.4]
  wire [1:0] _T_354; // @[Lookup.scala 11:37:@4246.4]
  wire [1:0] _T_355; // @[Lookup.scala 11:37:@4247.4]
  wire [1:0] _T_356; // @[Lookup.scala 11:37:@4248.4]
  wire [1:0] _T_357; // @[Lookup.scala 11:37:@4249.4]
  wire [2:0] _T_371; // @[Lookup.scala 11:37:@4264.4]
  wire [2:0] _T_372; // @[Lookup.scala 11:37:@4265.4]
  wire [2:0] _T_373; // @[Lookup.scala 11:37:@4266.4]
  wire [2:0] _T_374; // @[Lookup.scala 11:37:@4267.4]
  wire [2:0] _T_375; // @[Lookup.scala 11:37:@4268.4]
  wire [2:0] _T_376; // @[Lookup.scala 11:37:@4269.4]
  wire [2:0] _T_377; // @[Lookup.scala 11:37:@4270.4]
  wire [2:0] _T_378; // @[Lookup.scala 11:37:@4271.4]
  wire [2:0] _T_379; // @[Lookup.scala 11:37:@4272.4]
  wire [2:0] _T_380; // @[Lookup.scala 11:37:@4273.4]
  wire [2:0] _T_381; // @[Lookup.scala 11:37:@4274.4]
  wire [2:0] _T_382; // @[Lookup.scala 11:37:@4275.4]
  wire [2:0] _T_383; // @[Lookup.scala 11:37:@4276.4]
  wire [2:0] _T_384; // @[Lookup.scala 11:37:@4277.4]
  wire [2:0] _T_385; // @[Lookup.scala 11:37:@4278.4]
  wire [2:0] _T_386; // @[Lookup.scala 11:37:@4279.4]
  wire [2:0] _T_387; // @[Lookup.scala 11:37:@4280.4]
  wire [2:0] _T_388; // @[Lookup.scala 11:37:@4281.4]
  wire [2:0] _T_389; // @[Lookup.scala 11:37:@4282.4]
  wire [2:0] _T_390; // @[Lookup.scala 11:37:@4283.4]
  wire [2:0] _T_391; // @[Lookup.scala 11:37:@4284.4]
  wire [2:0] _T_392; // @[Lookup.scala 11:37:@4285.4]
  wire [2:0] _T_393; // @[Lookup.scala 11:37:@4286.4]
  wire [2:0] _T_394; // @[Lookup.scala 11:37:@4287.4]
  wire [2:0] _T_395; // @[Lookup.scala 11:37:@4288.4]
  wire [2:0] _T_396; // @[Lookup.scala 11:37:@4289.4]
  wire [2:0] _T_397; // @[Lookup.scala 11:37:@4290.4]
  wire [2:0] _T_398; // @[Lookup.scala 11:37:@4291.4]
  wire [2:0] _T_399; // @[Lookup.scala 11:37:@4292.4]
  wire [2:0] _T_400; // @[Lookup.scala 11:37:@4293.4]
  wire [2:0] _T_401; // @[Lookup.scala 11:37:@4294.4]
  wire [2:0] _T_402; // @[Lookup.scala 11:37:@4295.4]
  wire [2:0] _T_403; // @[Lookup.scala 11:37:@4296.4]
  wire [2:0] _T_404; // @[Lookup.scala 11:37:@4297.4]
  wire [2:0] _T_405; // @[Lookup.scala 11:37:@4298.4]
  wire [2:0] _T_406; // @[Lookup.scala 11:37:@4299.4]
  wire  _T_415; // @[Lookup.scala 11:37:@4309.4]
  wire  _T_416; // @[Lookup.scala 11:37:@4310.4]
  wire  _T_417; // @[Lookup.scala 11:37:@4311.4]
  wire  _T_418; // @[Lookup.scala 11:37:@4312.4]
  wire  _T_419; // @[Lookup.scala 11:37:@4313.4]
  wire  _T_420; // @[Lookup.scala 11:37:@4314.4]
  wire  _T_421; // @[Lookup.scala 11:37:@4315.4]
  wire  _T_422; // @[Lookup.scala 11:37:@4316.4]
  wire  _T_423; // @[Lookup.scala 11:37:@4317.4]
  wire  _T_424; // @[Lookup.scala 11:37:@4318.4]
  wire  _T_425; // @[Lookup.scala 11:37:@4319.4]
  wire  _T_426; // @[Lookup.scala 11:37:@4320.4]
  wire  _T_427; // @[Lookup.scala 11:37:@4321.4]
  wire  _T_428; // @[Lookup.scala 11:37:@4322.4]
  wire  _T_429; // @[Lookup.scala 11:37:@4323.4]
  wire  _T_430; // @[Lookup.scala 11:37:@4324.4]
  wire  _T_431; // @[Lookup.scala 11:37:@4325.4]
  wire  _T_432; // @[Lookup.scala 11:37:@4326.4]
  wire  _T_433; // @[Lookup.scala 11:37:@4327.4]
  wire  _T_434; // @[Lookup.scala 11:37:@4328.4]
  wire  _T_435; // @[Lookup.scala 11:37:@4329.4]
  wire  _T_436; // @[Lookup.scala 11:37:@4330.4]
  wire  _T_437; // @[Lookup.scala 11:37:@4331.4]
  wire  _T_438; // @[Lookup.scala 11:37:@4332.4]
  wire  _T_439; // @[Lookup.scala 11:37:@4333.4]
  wire  _T_440; // @[Lookup.scala 11:37:@4334.4]
  wire  _T_441; // @[Lookup.scala 11:37:@4335.4]
  wire  _T_442; // @[Lookup.scala 11:37:@4336.4]
  wire  _T_443; // @[Lookup.scala 11:37:@4337.4]
  wire  _T_444; // @[Lookup.scala 11:37:@4338.4]
  wire  _T_445; // @[Lookup.scala 11:37:@4339.4]
  wire  _T_446; // @[Lookup.scala 11:37:@4340.4]
  wire  _T_447; // @[Lookup.scala 11:37:@4341.4]
  wire  _T_448; // @[Lookup.scala 11:37:@4342.4]
  wire  _T_449; // @[Lookup.scala 11:37:@4343.4]
  wire  _T_450; // @[Lookup.scala 11:37:@4344.4]
  wire  _T_451; // @[Lookup.scala 11:37:@4345.4]
  wire  _T_452; // @[Lookup.scala 11:37:@4346.4]
  wire  _T_453; // @[Lookup.scala 11:37:@4347.4]
  wire  _T_454; // @[Lookup.scala 11:37:@4348.4]
  wire  _T_455; // @[Lookup.scala 11:37:@4349.4]
  wire  _T_475; // @[Lookup.scala 11:37:@4370.4]
  wire  _T_476; // @[Lookup.scala 11:37:@4371.4]
  wire  _T_477; // @[Lookup.scala 11:37:@4372.4]
  wire  _T_478; // @[Lookup.scala 11:37:@4373.4]
  wire  _T_479; // @[Lookup.scala 11:37:@4374.4]
  wire  _T_480; // @[Lookup.scala 11:37:@4375.4]
  wire  _T_481; // @[Lookup.scala 11:37:@4376.4]
  wire  _T_482; // @[Lookup.scala 11:37:@4377.4]
  wire  _T_483; // @[Lookup.scala 11:37:@4378.4]
  wire  _T_484; // @[Lookup.scala 11:37:@4379.4]
  wire  _T_485; // @[Lookup.scala 11:37:@4380.4]
  wire  _T_486; // @[Lookup.scala 11:37:@4381.4]
  wire  _T_487; // @[Lookup.scala 11:37:@4382.4]
  wire  _T_488; // @[Lookup.scala 11:37:@4383.4]
  wire  _T_489; // @[Lookup.scala 11:37:@4384.4]
  wire  _T_490; // @[Lookup.scala 11:37:@4385.4]
  wire  _T_491; // @[Lookup.scala 11:37:@4386.4]
  wire  _T_492; // @[Lookup.scala 11:37:@4387.4]
  wire  _T_493; // @[Lookup.scala 11:37:@4388.4]
  wire  _T_494; // @[Lookup.scala 11:37:@4389.4]
  wire  _T_495; // @[Lookup.scala 11:37:@4390.4]
  wire  _T_496; // @[Lookup.scala 11:37:@4391.4]
  wire  _T_497; // @[Lookup.scala 11:37:@4392.4]
  wire  _T_498; // @[Lookup.scala 11:37:@4393.4]
  wire  _T_499; // @[Lookup.scala 11:37:@4394.4]
  wire  _T_500; // @[Lookup.scala 11:37:@4395.4]
  wire  _T_501; // @[Lookup.scala 11:37:@4396.4]
  wire  _T_502; // @[Lookup.scala 11:37:@4397.4]
  wire  _T_503; // @[Lookup.scala 11:37:@4398.4]
  wire  _T_504; // @[Lookup.scala 11:37:@4399.4]
  wire [3:0] _T_512; // @[Lookup.scala 11:37:@4408.4]
  wire [3:0] _T_513; // @[Lookup.scala 11:37:@4409.4]
  wire [3:0] _T_514; // @[Lookup.scala 11:37:@4410.4]
  wire [3:0] _T_515; // @[Lookup.scala 11:37:@4411.4]
  wire [3:0] _T_516; // @[Lookup.scala 11:37:@4412.4]
  wire [3:0] _T_517; // @[Lookup.scala 11:37:@4413.4]
  wire [3:0] _T_518; // @[Lookup.scala 11:37:@4414.4]
  wire [3:0] _T_519; // @[Lookup.scala 11:37:@4415.4]
  wire [3:0] _T_520; // @[Lookup.scala 11:37:@4416.4]
  wire [3:0] _T_521; // @[Lookup.scala 11:37:@4417.4]
  wire [3:0] _T_522; // @[Lookup.scala 11:37:@4418.4]
  wire [3:0] _T_523; // @[Lookup.scala 11:37:@4419.4]
  wire [3:0] _T_524; // @[Lookup.scala 11:37:@4420.4]
  wire [3:0] _T_525; // @[Lookup.scala 11:37:@4421.4]
  wire [3:0] _T_526; // @[Lookup.scala 11:37:@4422.4]
  wire [3:0] _T_527; // @[Lookup.scala 11:37:@4423.4]
  wire [3:0] _T_528; // @[Lookup.scala 11:37:@4424.4]
  wire [3:0] _T_529; // @[Lookup.scala 11:37:@4425.4]
  wire [3:0] _T_530; // @[Lookup.scala 11:37:@4426.4]
  wire [3:0] _T_531; // @[Lookup.scala 11:37:@4427.4]
  wire [3:0] _T_532; // @[Lookup.scala 11:37:@4428.4]
  wire [3:0] _T_533; // @[Lookup.scala 11:37:@4429.4]
  wire [3:0] _T_534; // @[Lookup.scala 11:37:@4430.4]
  wire [3:0] _T_535; // @[Lookup.scala 11:37:@4431.4]
  wire [3:0] _T_536; // @[Lookup.scala 11:37:@4432.4]
  wire [3:0] _T_537; // @[Lookup.scala 11:37:@4433.4]
  wire [3:0] _T_538; // @[Lookup.scala 11:37:@4434.4]
  wire [3:0] _T_539; // @[Lookup.scala 11:37:@4435.4]
  wire [3:0] _T_540; // @[Lookup.scala 11:37:@4436.4]
  wire [3:0] _T_541; // @[Lookup.scala 11:37:@4437.4]
  wire [3:0] _T_542; // @[Lookup.scala 11:37:@4438.4]
  wire [3:0] _T_543; // @[Lookup.scala 11:37:@4439.4]
  wire [3:0] _T_544; // @[Lookup.scala 11:37:@4440.4]
  wire [3:0] _T_545; // @[Lookup.scala 11:37:@4441.4]
  wire [3:0] _T_546; // @[Lookup.scala 11:37:@4442.4]
  wire [3:0] _T_547; // @[Lookup.scala 11:37:@4443.4]
  wire [3:0] _T_548; // @[Lookup.scala 11:37:@4444.4]
  wire [3:0] _T_549; // @[Lookup.scala 11:37:@4445.4]
  wire [3:0] _T_550; // @[Lookup.scala 11:37:@4446.4]
  wire [3:0] _T_551; // @[Lookup.scala 11:37:@4447.4]
  wire [3:0] _T_552; // @[Lookup.scala 11:37:@4448.4]
  wire [3:0] _T_553; // @[Lookup.scala 11:37:@4449.4]
  wire [1:0] _T_561; // @[Lookup.scala 11:37:@4458.4]
  wire [1:0] _T_562; // @[Lookup.scala 11:37:@4459.4]
  wire [1:0] _T_563; // @[Lookup.scala 11:37:@4460.4]
  wire [1:0] _T_564; // @[Lookup.scala 11:37:@4461.4]
  wire [1:0] _T_565; // @[Lookup.scala 11:37:@4462.4]
  wire [1:0] _T_566; // @[Lookup.scala 11:37:@4463.4]
  wire [1:0] _T_567; // @[Lookup.scala 11:37:@4464.4]
  wire [1:0] _T_568; // @[Lookup.scala 11:37:@4465.4]
  wire [1:0] _T_569; // @[Lookup.scala 11:37:@4466.4]
  wire [1:0] _T_570; // @[Lookup.scala 11:37:@4467.4]
  wire [1:0] _T_571; // @[Lookup.scala 11:37:@4468.4]
  wire [1:0] _T_572; // @[Lookup.scala 11:37:@4469.4]
  wire [1:0] _T_573; // @[Lookup.scala 11:37:@4470.4]
  wire [1:0] _T_574; // @[Lookup.scala 11:37:@4471.4]
  wire [1:0] _T_575; // @[Lookup.scala 11:37:@4472.4]
  wire [1:0] _T_576; // @[Lookup.scala 11:37:@4473.4]
  wire [1:0] _T_577; // @[Lookup.scala 11:37:@4474.4]
  wire [1:0] _T_578; // @[Lookup.scala 11:37:@4475.4]
  wire [1:0] _T_579; // @[Lookup.scala 11:37:@4476.4]
  wire [1:0] _T_580; // @[Lookup.scala 11:37:@4477.4]
  wire [1:0] _T_581; // @[Lookup.scala 11:37:@4478.4]
  wire [1:0] _T_582; // @[Lookup.scala 11:37:@4479.4]
  wire [1:0] _T_583; // @[Lookup.scala 11:37:@4480.4]
  wire [1:0] _T_584; // @[Lookup.scala 11:37:@4481.4]
  wire [1:0] _T_585; // @[Lookup.scala 11:37:@4482.4]
  wire [1:0] _T_586; // @[Lookup.scala 11:37:@4483.4]
  wire [1:0] _T_587; // @[Lookup.scala 11:37:@4484.4]
  wire [1:0] _T_588; // @[Lookup.scala 11:37:@4485.4]
  wire [1:0] _T_589; // @[Lookup.scala 11:37:@4486.4]
  wire [1:0] _T_590; // @[Lookup.scala 11:37:@4487.4]
  wire [1:0] _T_591; // @[Lookup.scala 11:37:@4488.4]
  wire [1:0] _T_592; // @[Lookup.scala 11:37:@4489.4]
  wire [1:0] _T_593; // @[Lookup.scala 11:37:@4490.4]
  wire [1:0] _T_594; // @[Lookup.scala 11:37:@4491.4]
  wire [1:0] _T_595; // @[Lookup.scala 11:37:@4492.4]
  wire [1:0] _T_596; // @[Lookup.scala 11:37:@4493.4]
  wire [1:0] _T_597; // @[Lookup.scala 11:37:@4494.4]
  wire [1:0] _T_598; // @[Lookup.scala 11:37:@4495.4]
  wire [1:0] _T_599; // @[Lookup.scala 11:37:@4496.4]
  wire [1:0] _T_600; // @[Lookup.scala 11:37:@4497.4]
  wire [1:0] _T_601; // @[Lookup.scala 11:37:@4498.4]
  wire [1:0] _T_602; // @[Lookup.scala 11:37:@4499.4]
  wire  _T_616; // @[Lookup.scala 11:37:@4514.4]
  wire  _T_617; // @[Lookup.scala 11:37:@4515.4]
  wire  _T_618; // @[Lookup.scala 11:37:@4516.4]
  wire  _T_619; // @[Lookup.scala 11:37:@4517.4]
  wire  _T_620; // @[Lookup.scala 11:37:@4518.4]
  wire  _T_621; // @[Lookup.scala 11:37:@4519.4]
  wire  _T_622; // @[Lookup.scala 11:37:@4520.4]
  wire  _T_623; // @[Lookup.scala 11:37:@4521.4]
  wire  _T_624; // @[Lookup.scala 11:37:@4522.4]
  wire  _T_625; // @[Lookup.scala 11:37:@4523.4]
  wire  _T_626; // @[Lookup.scala 11:37:@4524.4]
  wire  _T_627; // @[Lookup.scala 11:37:@4525.4]
  wire  _T_628; // @[Lookup.scala 11:37:@4526.4]
  wire  _T_629; // @[Lookup.scala 11:37:@4527.4]
  wire  _T_630; // @[Lookup.scala 11:37:@4528.4]
  wire  _T_631; // @[Lookup.scala 11:37:@4529.4]
  wire  _T_632; // @[Lookup.scala 11:37:@4530.4]
  wire  _T_633; // @[Lookup.scala 11:37:@4531.4]
  wire  _T_634; // @[Lookup.scala 11:37:@4532.4]
  wire  _T_635; // @[Lookup.scala 11:37:@4533.4]
  wire  _T_636; // @[Lookup.scala 11:37:@4534.4]
  wire  _T_637; // @[Lookup.scala 11:37:@4535.4]
  wire  _T_638; // @[Lookup.scala 11:37:@4536.4]
  wire  _T_639; // @[Lookup.scala 11:37:@4537.4]
  wire  _T_640; // @[Lookup.scala 11:37:@4538.4]
  wire  _T_641; // @[Lookup.scala 11:37:@4539.4]
  wire  _T_642; // @[Lookup.scala 11:37:@4540.4]
  wire  _T_643; // @[Lookup.scala 11:37:@4541.4]
  wire  _T_644; // @[Lookup.scala 11:37:@4542.4]
  wire  _T_645; // @[Lookup.scala 11:37:@4543.4]
  wire  _T_646; // @[Lookup.scala 11:37:@4544.4]
  wire  _T_647; // @[Lookup.scala 11:37:@4545.4]
  wire  _T_648; // @[Lookup.scala 11:37:@4546.4]
  wire  _T_649; // @[Lookup.scala 11:37:@4547.4]
  wire  _T_650; // @[Lookup.scala 11:37:@4548.4]
  wire  _T_651; // @[Lookup.scala 11:37:@4549.4]
  wire  _T_653; // @[Lookup.scala 11:37:@4552.4]
  wire  _T_654; // @[Lookup.scala 11:37:@4553.4]
  wire  _T_655; // @[Lookup.scala 11:37:@4554.4]
  wire  _T_656; // @[Lookup.scala 11:37:@4555.4]
  wire  _T_657; // @[Lookup.scala 11:37:@4556.4]
  wire  _T_658; // @[Lookup.scala 11:37:@4557.4]
  wire  _T_659; // @[Lookup.scala 11:37:@4558.4]
  wire  _T_660; // @[Lookup.scala 11:37:@4559.4]
  wire  _T_661; // @[Lookup.scala 11:37:@4560.4]
  wire  _T_662; // @[Lookup.scala 11:37:@4561.4]
  wire  _T_663; // @[Lookup.scala 11:37:@4562.4]
  wire  _T_664; // @[Lookup.scala 11:37:@4563.4]
  wire  _T_665; // @[Lookup.scala 11:37:@4564.4]
  wire  _T_666; // @[Lookup.scala 11:37:@4565.4]
  wire  _T_667; // @[Lookup.scala 11:37:@4566.4]
  wire  _T_668; // @[Lookup.scala 11:37:@4567.4]
  wire  _T_669; // @[Lookup.scala 11:37:@4568.4]
  wire  _T_670; // @[Lookup.scala 11:37:@4569.4]
  wire  _T_671; // @[Lookup.scala 11:37:@4570.4]
  wire  _T_672; // @[Lookup.scala 11:37:@4571.4]
  wire  _T_673; // @[Lookup.scala 11:37:@4572.4]
  wire  _T_674; // @[Lookup.scala 11:37:@4573.4]
  wire  _T_675; // @[Lookup.scala 11:37:@4574.4]
  wire  _T_676; // @[Lookup.scala 11:37:@4575.4]
  wire  _T_677; // @[Lookup.scala 11:37:@4576.4]
  wire  _T_678; // @[Lookup.scala 11:37:@4577.4]
  wire  _T_679; // @[Lookup.scala 11:37:@4578.4]
  wire  _T_680; // @[Lookup.scala 11:37:@4579.4]
  wire  _T_681; // @[Lookup.scala 11:37:@4580.4]
  wire  _T_682; // @[Lookup.scala 11:37:@4581.4]
  wire  _T_683; // @[Lookup.scala 11:37:@4582.4]
  wire  _T_684; // @[Lookup.scala 11:37:@4583.4]
  wire  _T_685; // @[Lookup.scala 11:37:@4584.4]
  wire  _T_686; // @[Lookup.scala 11:37:@4585.4]
  wire  _T_687; // @[Lookup.scala 11:37:@4586.4]
  wire  _T_688; // @[Lookup.scala 11:37:@4587.4]
  wire  _T_689; // @[Lookup.scala 11:37:@4588.4]
  wire  _T_690; // @[Lookup.scala 11:37:@4589.4]
  wire  _T_691; // @[Lookup.scala 11:37:@4590.4]
  wire  _T_692; // @[Lookup.scala 11:37:@4591.4]
  wire  _T_693; // @[Lookup.scala 11:37:@4592.4]
  wire  _T_694; // @[Lookup.scala 11:37:@4593.4]
  wire  _T_695; // @[Lookup.scala 11:37:@4594.4]
  wire  _T_696; // @[Lookup.scala 11:37:@4595.4]
  wire  _T_697; // @[Lookup.scala 11:37:@4596.4]
  wire  _T_698; // @[Lookup.scala 11:37:@4597.4]
  wire  _T_699; // @[Lookup.scala 11:37:@4598.4]
  wire  _T_700; // @[Lookup.scala 11:37:@4599.4]
  wire  _T_744; // @[Lookup.scala 11:37:@4644.4]
  wire  _T_745; // @[Lookup.scala 11:37:@4645.4]
  wire  _T_746; // @[Lookup.scala 11:37:@4646.4]
  wire  _T_747; // @[Lookup.scala 11:37:@4647.4]
  wire  _T_748; // @[Lookup.scala 11:37:@4648.4]
  wire  _T_749; // @[Lookup.scala 11:37:@4649.4]
  wire [2:0] _T_792; // @[Lookup.scala 11:37:@4693.4]
  wire [2:0] _T_793; // @[Lookup.scala 11:37:@4694.4]
  wire [2:0] _T_794; // @[Lookup.scala 11:37:@4695.4]
  wire [2:0] _T_795; // @[Lookup.scala 11:37:@4696.4]
  wire [2:0] _T_796; // @[Lookup.scala 11:37:@4697.4]
  wire [2:0] _T_797; // @[Lookup.scala 11:37:@4698.4]
  wire [2:0] _T_798; // @[Lookup.scala 11:37:@4699.4]
  wire [2:0] _T_802; // @[Lookup.scala 11:37:@4704.4]
  wire [2:0] _T_803; // @[Lookup.scala 11:37:@4705.4]
  wire [2:0] _T_804; // @[Lookup.scala 11:37:@4706.4]
  wire [2:0] _T_805; // @[Lookup.scala 11:37:@4707.4]
  wire [2:0] _T_806; // @[Lookup.scala 11:37:@4708.4]
  wire [2:0] _T_807; // @[Lookup.scala 11:37:@4709.4]
  wire [2:0] _T_808; // @[Lookup.scala 11:37:@4710.4]
  wire [2:0] _T_809; // @[Lookup.scala 11:37:@4711.4]
  wire [2:0] _T_810; // @[Lookup.scala 11:37:@4712.4]
  wire [2:0] _T_811; // @[Lookup.scala 11:37:@4713.4]
  wire [2:0] _T_812; // @[Lookup.scala 11:37:@4714.4]
  wire [2:0] _T_813; // @[Lookup.scala 11:37:@4715.4]
  wire [2:0] _T_814; // @[Lookup.scala 11:37:@4716.4]
  wire [2:0] _T_815; // @[Lookup.scala 11:37:@4717.4]
  wire [2:0] _T_816; // @[Lookup.scala 11:37:@4718.4]
  wire [2:0] _T_817; // @[Lookup.scala 11:37:@4719.4]
  wire [2:0] _T_818; // @[Lookup.scala 11:37:@4720.4]
  wire [2:0] _T_819; // @[Lookup.scala 11:37:@4721.4]
  wire [2:0] _T_820; // @[Lookup.scala 11:37:@4722.4]
  wire [2:0] _T_821; // @[Lookup.scala 11:37:@4723.4]
  wire [2:0] _T_822; // @[Lookup.scala 11:37:@4724.4]
  wire [2:0] _T_823; // @[Lookup.scala 11:37:@4725.4]
  wire [2:0] _T_824; // @[Lookup.scala 11:37:@4726.4]
  wire [2:0] _T_825; // @[Lookup.scala 11:37:@4727.4]
  wire [2:0] _T_826; // @[Lookup.scala 11:37:@4728.4]
  wire [2:0] _T_827; // @[Lookup.scala 11:37:@4729.4]
  wire [2:0] _T_828; // @[Lookup.scala 11:37:@4730.4]
  wire [2:0] _T_829; // @[Lookup.scala 11:37:@4731.4]
  wire [2:0] _T_830; // @[Lookup.scala 11:37:@4732.4]
  wire [2:0] _T_831; // @[Lookup.scala 11:37:@4733.4]
  wire [2:0] _T_832; // @[Lookup.scala 11:37:@4734.4]
  wire [2:0] _T_833; // @[Lookup.scala 11:37:@4735.4]
  wire [2:0] _T_834; // @[Lookup.scala 11:37:@4736.4]
  wire [2:0] _T_835; // @[Lookup.scala 11:37:@4737.4]
  wire [2:0] _T_836; // @[Lookup.scala 11:37:@4738.4]
  wire [2:0] _T_837; // @[Lookup.scala 11:37:@4739.4]
  wire [2:0] _T_838; // @[Lookup.scala 11:37:@4740.4]
  wire [2:0] _T_839; // @[Lookup.scala 11:37:@4741.4]
  wire [2:0] _T_840; // @[Lookup.scala 11:37:@4742.4]
  wire [2:0] _T_841; // @[Lookup.scala 11:37:@4743.4]
  wire [2:0] _T_842; // @[Lookup.scala 11:37:@4744.4]
  wire [2:0] _T_843; // @[Lookup.scala 11:37:@4745.4]
  wire [2:0] _T_844; // @[Lookup.scala 11:37:@4746.4]
  wire [2:0] _T_845; // @[Lookup.scala 11:37:@4747.4]
  wire [2:0] _T_846; // @[Lookup.scala 11:37:@4748.4]
  wire [2:0] _T_847; // @[Lookup.scala 11:37:@4749.4]
  wire  _T_850; // @[Lookup.scala 11:37:@4753.4]
  wire  _T_851; // @[Lookup.scala 11:37:@4754.4]
  wire  _T_852; // @[Lookup.scala 11:37:@4755.4]
  wire  _T_853; // @[Lookup.scala 11:37:@4756.4]
  wire  _T_854; // @[Lookup.scala 11:37:@4757.4]
  wire  _T_855; // @[Lookup.scala 11:37:@4758.4]
  wire  _T_856; // @[Lookup.scala 11:37:@4759.4]
  wire  _T_857; // @[Lookup.scala 11:37:@4760.4]
  wire  _T_858; // @[Lookup.scala 11:37:@4761.4]
  wire  _T_859; // @[Lookup.scala 11:37:@4762.4]
  wire  _T_860; // @[Lookup.scala 11:37:@4763.4]
  wire  _T_861; // @[Lookup.scala 11:37:@4764.4]
  wire  _T_862; // @[Lookup.scala 11:37:@4765.4]
  wire  _T_863; // @[Lookup.scala 11:37:@4766.4]
  wire  _T_864; // @[Lookup.scala 11:37:@4767.4]
  wire  _T_865; // @[Lookup.scala 11:37:@4768.4]
  wire  _T_866; // @[Lookup.scala 11:37:@4769.4]
  wire  _T_867; // @[Lookup.scala 11:37:@4770.4]
  wire  _T_868; // @[Lookup.scala 11:37:@4771.4]
  wire  _T_869; // @[Lookup.scala 11:37:@4772.4]
  wire  _T_870; // @[Lookup.scala 11:37:@4773.4]
  wire  _T_871; // @[Lookup.scala 11:37:@4774.4]
  wire  _T_872; // @[Lookup.scala 11:37:@4775.4]
  wire  _T_873; // @[Lookup.scala 11:37:@4776.4]
  wire  _T_874; // @[Lookup.scala 11:37:@4777.4]
  wire  _T_875; // @[Lookup.scala 11:37:@4778.4]
  wire  _T_876; // @[Lookup.scala 11:37:@4779.4]
  wire  _T_877; // @[Lookup.scala 11:37:@4780.4]
  wire  _T_878; // @[Lookup.scala 11:37:@4781.4]
  wire  _T_879; // @[Lookup.scala 11:37:@4782.4]
  wire  _T_880; // @[Lookup.scala 11:37:@4783.4]
  wire  _T_881; // @[Lookup.scala 11:37:@4784.4]
  wire  _T_882; // @[Lookup.scala 11:37:@4785.4]
  wire  _T_883; // @[Lookup.scala 11:37:@4786.4]
  wire  _T_884; // @[Lookup.scala 11:37:@4787.4]
  wire  _T_885; // @[Lookup.scala 11:37:@4788.4]
  wire  _T_886; // @[Lookup.scala 11:37:@4789.4]
  wire  _T_887; // @[Lookup.scala 11:37:@4790.4]
  wire  _T_888; // @[Lookup.scala 11:37:@4791.4]
  wire  _T_889; // @[Lookup.scala 11:37:@4792.4]
  wire  _T_890; // @[Lookup.scala 11:37:@4793.4]
  wire  _T_891; // @[Lookup.scala 11:37:@4794.4]
  wire  _T_892; // @[Lookup.scala 11:37:@4795.4]
  wire  _T_893; // @[Lookup.scala 11:37:@4796.4]
  wire  _T_894; // @[Lookup.scala 11:37:@4797.4]
  wire  _T_895; // @[Lookup.scala 11:37:@4798.4]
  wire  _T_896; // @[Lookup.scala 11:37:@4799.4]
  wire [4:0] _T_899; // @[InstDecoder.scala 130:31:@4816.4]
  wire [4:0] _T_901; // @[InstDecoder.scala 132:31:@4820.4]
  wire [4:0] func; // @[InstDecoder.scala 134:21:@4822.4]
  wire  _T_905; // @[InstDecoder.scala 136:38:@4825.4]
  wire  _T_907; // @[InstDecoder.scala 137:39:@4826.4]
  wire  _T_908; // @[InstDecoder.scala 141:32:@4827.4]
  wire  _T_910; // @[InstDecoder.scala 135:37:@4828.4]
  wire  _T_912; // @[InstDecoder.scala 135:53:@4829.4]
  wire  _T_913; // @[InstDecoder.scala 135:45:@4830.4]
  wire [4:0] _GEN_0; // @[InstDecoder.scala 142:24:@4834.4]
  wire  _T_917; // @[InstDecoder.scala 142:24:@4834.4]
  wire  _T_919; // @[InstDecoder.scala 135:37:@4835.4]
  wire  _T_921; // @[InstDecoder.scala 135:53:@4836.4]
  wire  _T_922; // @[InstDecoder.scala 135:45:@4837.4]
  wire  _T_923; // @[InstDecoder.scala 142:41:@4838.4]
  wire  _T_930; // @[InstDecoder.scala 143:6:@4842.4]
  wire  _T_931; // @[InstDecoder.scala 143:50:@4843.4]
  wire  _T_932; // @[InstDecoder.scala 143:29:@4844.4]
  wire [11:0] imm_itype; // @[InstDecoder.scala 146:27:@4847.4]
  wire [6:0] _T_934; // @[InstDecoder.scala 147:31:@4848.4]
  wire [11:0] imm_stype; // @[Cat.scala 30:58:@4850.4]
  wire  _T_936; // @[InstDecoder.scala 148:31:@4851.4]
  wire  _T_937; // @[InstDecoder.scala 148:44:@4852.4]
  wire [5:0] _T_938; // @[InstDecoder.scala 148:56:@4853.4]
  wire [3:0] _T_939; // @[InstDecoder.scala 148:73:@4854.4]
  wire [11:0] imm_sbtype; // @[Cat.scala 30:58:@4857.4]
  wire [19:0] imm_utype; // @[InstDecoder.scala 149:27:@4858.4]
  wire [7:0] _T_943; // @[InstDecoder.scala 150:44:@4860.4]
  wire  _T_944; // @[InstDecoder.scala 150:60:@4861.4]
  wire [9:0] _T_945; // @[InstDecoder.scala 150:73:@4862.4]
  wire [19:0] imm_ujtype; // @[Cat.scala 30:58:@4865.4]
  wire  _T_948; // @[InstDecoder.scala 153:43:@4866.4]
  wire [19:0] _T_952; // @[Bitwise.scala 72:12:@4868.4]
  wire  _T_954; // @[InstDecoder.scala 154:43:@4871.4]
  wire [19:0] _T_958; // @[Bitwise.scala 72:12:@4873.4]
  wire  _T_960; // @[InstDecoder.scala 155:44:@4876.4]
  wire [18:0] _T_964; // @[Bitwise.scala 72:12:@4878.4]
  wire [30:0] _T_966; // @[Cat.scala 30:58:@4879.4]
  wire  _T_974; // @[InstDecoder.scala 157:44:@4885.4]
  wire [10:0] _T_978; // @[Bitwise.scala 72:12:@4887.4]
  wire [30:0] _T_980; // @[Cat.scala 30:58:@4888.4]
  assign _T_13 = io_inst & 32'h707f; // @[Lookup.scala 9:38:@4001.4]
  assign _T_14 = 32'h2003 == _T_13; // @[Lookup.scala 9:38:@4002.4]
  assign _T_18 = 32'h3 == _T_13; // @[Lookup.scala 9:38:@4004.4]
  assign _T_22 = 32'h4003 == _T_13; // @[Lookup.scala 9:38:@4006.4]
  assign _T_26 = 32'h1003 == _T_13; // @[Lookup.scala 9:38:@4008.4]
  assign _T_30 = 32'h5003 == _T_13; // @[Lookup.scala 9:38:@4010.4]
  assign _T_34 = 32'h2023 == _T_13; // @[Lookup.scala 9:38:@4012.4]
  assign _T_38 = 32'h23 == _T_13; // @[Lookup.scala 9:38:@4014.4]
  assign _T_42 = 32'h1023 == _T_13; // @[Lookup.scala 9:38:@4016.4]
  assign _T_45 = io_inst & 32'h7f; // @[Lookup.scala 9:38:@4017.4]
  assign _T_46 = 32'h17 == _T_45; // @[Lookup.scala 9:38:@4018.4]
  assign _T_50 = 32'h37 == _T_45; // @[Lookup.scala 9:38:@4020.4]
  assign _T_54 = 32'h13 == _T_13; // @[Lookup.scala 9:38:@4022.4]
  assign _T_58 = 32'h7013 == _T_13; // @[Lookup.scala 9:38:@4024.4]
  assign _T_62 = 32'h6013 == _T_13; // @[Lookup.scala 9:38:@4026.4]
  assign _T_66 = 32'h4013 == _T_13; // @[Lookup.scala 9:38:@4028.4]
  assign _T_70 = 32'h2013 == _T_13; // @[Lookup.scala 9:38:@4030.4]
  assign _T_74 = 32'h3013 == _T_13; // @[Lookup.scala 9:38:@4032.4]
  assign _T_77 = io_inst & 32'hfc00707f; // @[Lookup.scala 9:38:@4033.4]
  assign _T_78 = 32'h1013 == _T_77; // @[Lookup.scala 9:38:@4034.4]
  assign _T_82 = 32'h40005013 == _T_77; // @[Lookup.scala 9:38:@4036.4]
  assign _T_86 = 32'h5013 == _T_77; // @[Lookup.scala 9:38:@4038.4]
  assign _T_89 = io_inst & 32'hfe00707f; // @[Lookup.scala 9:38:@4039.4]
  assign _T_90 = 32'h1033 == _T_89; // @[Lookup.scala 9:38:@4040.4]
  assign _T_94 = 32'h33 == _T_89; // @[Lookup.scala 9:38:@4042.4]
  assign _T_98 = 32'h40000033 == _T_89; // @[Lookup.scala 9:38:@4044.4]
  assign _T_102 = 32'h2033 == _T_89; // @[Lookup.scala 9:38:@4046.4]
  assign _T_106 = 32'h3033 == _T_89; // @[Lookup.scala 9:38:@4048.4]
  assign _T_110 = 32'h7033 == _T_89; // @[Lookup.scala 9:38:@4050.4]
  assign _T_114 = 32'h6033 == _T_89; // @[Lookup.scala 9:38:@4052.4]
  assign _T_118 = 32'h4033 == _T_89; // @[Lookup.scala 9:38:@4054.4]
  assign _T_122 = 32'h40005033 == _T_89; // @[Lookup.scala 9:38:@4056.4]
  assign _T_126 = 32'h5033 == _T_89; // @[Lookup.scala 9:38:@4058.4]
  assign _T_130 = 32'h6f == _T_45; // @[Lookup.scala 9:38:@4060.4]
  assign _T_134 = 32'h67 == _T_13; // @[Lookup.scala 9:38:@4062.4]
  assign _T_138 = 32'h63 == _T_13; // @[Lookup.scala 9:38:@4064.4]
  assign _T_142 = 32'h1063 == _T_13; // @[Lookup.scala 9:38:@4066.4]
  assign _T_146 = 32'h5063 == _T_13; // @[Lookup.scala 9:38:@4068.4]
  assign _T_150 = 32'h7063 == _T_13; // @[Lookup.scala 9:38:@4070.4]
  assign _T_154 = 32'h4063 == _T_13; // @[Lookup.scala 9:38:@4072.4]
  assign _T_158 = 32'h6063 == _T_13; // @[Lookup.scala 9:38:@4074.4]
  assign _T_162 = 32'h5073 == _T_13; // @[Lookup.scala 9:38:@4076.4]
  assign _T_166 = 32'h6073 == _T_13; // @[Lookup.scala 9:38:@4078.4]
  assign _T_170 = 32'h1073 == _T_13; // @[Lookup.scala 9:38:@4080.4]
  assign _T_174 = 32'h2073 == _T_13; // @[Lookup.scala 9:38:@4082.4]
  assign _T_178 = 32'h3073 == _T_13; // @[Lookup.scala 9:38:@4084.4]
  assign _T_182 = 32'h7073 == _T_13; // @[Lookup.scala 9:38:@4086.4]
  assign _T_186 = 32'h73 == io_inst; // @[Lookup.scala 9:38:@4088.4]
  assign _T_190 = 32'h30200073 == io_inst; // @[Lookup.scala 9:38:@4090.4]
  assign _T_194 = 32'h7b200073 == io_inst; // @[Lookup.scala 9:38:@4092.4]
  assign _T_198 = 32'h100073 == io_inst; // @[Lookup.scala 9:38:@4094.4]
  assign _T_202 = 32'h10500073 == io_inst; // @[Lookup.scala 9:38:@4096.4]
  assign _T_206 = 32'h100f == _T_13; // @[Lookup.scala 9:38:@4098.4]
  assign _T_210 = 32'hf == _T_13; // @[Lookup.scala 9:38:@4100.4]
  assign _T_212 = _T_206 ? 1'h1 : _T_210; // @[Lookup.scala 11:37:@4102.4]
  assign _T_213 = _T_202 ? 1'h1 : _T_212; // @[Lookup.scala 11:37:@4103.4]
  assign _T_214 = _T_198 ? 1'h1 : _T_213; // @[Lookup.scala 11:37:@4104.4]
  assign _T_215 = _T_194 ? 1'h1 : _T_214; // @[Lookup.scala 11:37:@4105.4]
  assign _T_216 = _T_190 ? 1'h1 : _T_215; // @[Lookup.scala 11:37:@4106.4]
  assign _T_217 = _T_186 ? 1'h1 : _T_216; // @[Lookup.scala 11:37:@4107.4]
  assign _T_218 = _T_182 ? 1'h1 : _T_217; // @[Lookup.scala 11:37:@4108.4]
  assign _T_219 = _T_178 ? 1'h1 : _T_218; // @[Lookup.scala 11:37:@4109.4]
  assign _T_220 = _T_174 ? 1'h1 : _T_219; // @[Lookup.scala 11:37:@4110.4]
  assign _T_221 = _T_170 ? 1'h1 : _T_220; // @[Lookup.scala 11:37:@4111.4]
  assign _T_222 = _T_166 ? 1'h1 : _T_221; // @[Lookup.scala 11:37:@4112.4]
  assign _T_223 = _T_162 ? 1'h1 : _T_222; // @[Lookup.scala 11:37:@4113.4]
  assign _T_224 = _T_158 ? 1'h1 : _T_223; // @[Lookup.scala 11:37:@4114.4]
  assign _T_225 = _T_154 ? 1'h1 : _T_224; // @[Lookup.scala 11:37:@4115.4]
  assign _T_226 = _T_150 ? 1'h1 : _T_225; // @[Lookup.scala 11:37:@4116.4]
  assign _T_227 = _T_146 ? 1'h1 : _T_226; // @[Lookup.scala 11:37:@4117.4]
  assign _T_228 = _T_142 ? 1'h1 : _T_227; // @[Lookup.scala 11:37:@4118.4]
  assign _T_229 = _T_138 ? 1'h1 : _T_228; // @[Lookup.scala 11:37:@4119.4]
  assign _T_230 = _T_134 ? 1'h1 : _T_229; // @[Lookup.scala 11:37:@4120.4]
  assign _T_231 = _T_130 ? 1'h1 : _T_230; // @[Lookup.scala 11:37:@4121.4]
  assign _T_232 = _T_126 ? 1'h1 : _T_231; // @[Lookup.scala 11:37:@4122.4]
  assign _T_233 = _T_122 ? 1'h1 : _T_232; // @[Lookup.scala 11:37:@4123.4]
  assign _T_234 = _T_118 ? 1'h1 : _T_233; // @[Lookup.scala 11:37:@4124.4]
  assign _T_235 = _T_114 ? 1'h1 : _T_234; // @[Lookup.scala 11:37:@4125.4]
  assign _T_236 = _T_110 ? 1'h1 : _T_235; // @[Lookup.scala 11:37:@4126.4]
  assign _T_237 = _T_106 ? 1'h1 : _T_236; // @[Lookup.scala 11:37:@4127.4]
  assign _T_238 = _T_102 ? 1'h1 : _T_237; // @[Lookup.scala 11:37:@4128.4]
  assign _T_239 = _T_98 ? 1'h1 : _T_238; // @[Lookup.scala 11:37:@4129.4]
  assign _T_240 = _T_94 ? 1'h1 : _T_239; // @[Lookup.scala 11:37:@4130.4]
  assign _T_241 = _T_90 ? 1'h1 : _T_240; // @[Lookup.scala 11:37:@4131.4]
  assign _T_242 = _T_86 ? 1'h1 : _T_241; // @[Lookup.scala 11:37:@4132.4]
  assign _T_243 = _T_82 ? 1'h1 : _T_242; // @[Lookup.scala 11:37:@4133.4]
  assign _T_244 = _T_78 ? 1'h1 : _T_243; // @[Lookup.scala 11:37:@4134.4]
  assign _T_245 = _T_74 ? 1'h1 : _T_244; // @[Lookup.scala 11:37:@4135.4]
  assign _T_246 = _T_70 ? 1'h1 : _T_245; // @[Lookup.scala 11:37:@4136.4]
  assign _T_247 = _T_66 ? 1'h1 : _T_246; // @[Lookup.scala 11:37:@4137.4]
  assign _T_248 = _T_62 ? 1'h1 : _T_247; // @[Lookup.scala 11:37:@4138.4]
  assign _T_249 = _T_58 ? 1'h1 : _T_248; // @[Lookup.scala 11:37:@4139.4]
  assign _T_250 = _T_54 ? 1'h1 : _T_249; // @[Lookup.scala 11:37:@4140.4]
  assign _T_251 = _T_50 ? 1'h1 : _T_250; // @[Lookup.scala 11:37:@4141.4]
  assign _T_252 = _T_46 ? 1'h1 : _T_251; // @[Lookup.scala 11:37:@4142.4]
  assign _T_253 = _T_42 ? 1'h1 : _T_252; // @[Lookup.scala 11:37:@4143.4]
  assign _T_254 = _T_38 ? 1'h1 : _T_253; // @[Lookup.scala 11:37:@4144.4]
  assign _T_255 = _T_34 ? 1'h1 : _T_254; // @[Lookup.scala 11:37:@4145.4]
  assign _T_256 = _T_30 ? 1'h1 : _T_255; // @[Lookup.scala 11:37:@4146.4]
  assign _T_257 = _T_26 ? 1'h1 : _T_256; // @[Lookup.scala 11:37:@4147.4]
  assign _T_258 = _T_22 ? 1'h1 : _T_257; // @[Lookup.scala 11:37:@4148.4]
  assign _T_259 = _T_18 ? 1'h1 : _T_258; // @[Lookup.scala 11:37:@4149.4]
  assign signals_0 = _T_14 ? 1'h1 : _T_259; // @[Lookup.scala 11:37:@4150.4]
  assign _T_273 = _T_158 ? 4'h6 : 4'h0; // @[Lookup.scala 11:37:@4164.4]
  assign _T_274 = _T_154 ? 4'h5 : _T_273; // @[Lookup.scala 11:37:@4165.4]
  assign _T_275 = _T_150 ? 4'h4 : _T_274; // @[Lookup.scala 11:37:@4166.4]
  assign _T_276 = _T_146 ? 4'h3 : _T_275; // @[Lookup.scala 11:37:@4167.4]
  assign _T_277 = _T_142 ? 4'h1 : _T_276; // @[Lookup.scala 11:37:@4168.4]
  assign _T_278 = _T_138 ? 4'h2 : _T_277; // @[Lookup.scala 11:37:@4169.4]
  assign _T_279 = _T_134 ? 4'h8 : _T_278; // @[Lookup.scala 11:37:@4170.4]
  assign _T_280 = _T_130 ? 4'h7 : _T_279; // @[Lookup.scala 11:37:@4171.4]
  assign _T_281 = _T_126 ? 4'h0 : _T_280; // @[Lookup.scala 11:37:@4172.4]
  assign _T_282 = _T_122 ? 4'h0 : _T_281; // @[Lookup.scala 11:37:@4173.4]
  assign _T_283 = _T_118 ? 4'h0 : _T_282; // @[Lookup.scala 11:37:@4174.4]
  assign _T_284 = _T_114 ? 4'h0 : _T_283; // @[Lookup.scala 11:37:@4175.4]
  assign _T_285 = _T_110 ? 4'h0 : _T_284; // @[Lookup.scala 11:37:@4176.4]
  assign _T_286 = _T_106 ? 4'h0 : _T_285; // @[Lookup.scala 11:37:@4177.4]
  assign _T_287 = _T_102 ? 4'h0 : _T_286; // @[Lookup.scala 11:37:@4178.4]
  assign _T_288 = _T_98 ? 4'h0 : _T_287; // @[Lookup.scala 11:37:@4179.4]
  assign _T_289 = _T_94 ? 4'h0 : _T_288; // @[Lookup.scala 11:37:@4180.4]
  assign _T_290 = _T_90 ? 4'h0 : _T_289; // @[Lookup.scala 11:37:@4181.4]
  assign _T_291 = _T_86 ? 4'h0 : _T_290; // @[Lookup.scala 11:37:@4182.4]
  assign _T_292 = _T_82 ? 4'h0 : _T_291; // @[Lookup.scala 11:37:@4183.4]
  assign _T_293 = _T_78 ? 4'h0 : _T_292; // @[Lookup.scala 11:37:@4184.4]
  assign _T_294 = _T_74 ? 4'h0 : _T_293; // @[Lookup.scala 11:37:@4185.4]
  assign _T_295 = _T_70 ? 4'h0 : _T_294; // @[Lookup.scala 11:37:@4186.4]
  assign _T_296 = _T_66 ? 4'h0 : _T_295; // @[Lookup.scala 11:37:@4187.4]
  assign _T_297 = _T_62 ? 4'h0 : _T_296; // @[Lookup.scala 11:37:@4188.4]
  assign _T_298 = _T_58 ? 4'h0 : _T_297; // @[Lookup.scala 11:37:@4189.4]
  assign _T_299 = _T_54 ? 4'h0 : _T_298; // @[Lookup.scala 11:37:@4190.4]
  assign _T_300 = _T_50 ? 4'h0 : _T_299; // @[Lookup.scala 11:37:@4191.4]
  assign _T_301 = _T_46 ? 4'h0 : _T_300; // @[Lookup.scala 11:37:@4192.4]
  assign _T_302 = _T_42 ? 4'h0 : _T_301; // @[Lookup.scala 11:37:@4193.4]
  assign _T_303 = _T_38 ? 4'h0 : _T_302; // @[Lookup.scala 11:37:@4194.4]
  assign _T_304 = _T_34 ? 4'h0 : _T_303; // @[Lookup.scala 11:37:@4195.4]
  assign _T_305 = _T_30 ? 4'h0 : _T_304; // @[Lookup.scala 11:37:@4196.4]
  assign _T_306 = _T_26 ? 4'h0 : _T_305; // @[Lookup.scala 11:37:@4197.4]
  assign _T_307 = _T_22 ? 4'h0 : _T_306; // @[Lookup.scala 11:37:@4198.4]
  assign _T_308 = _T_18 ? 4'h0 : _T_307; // @[Lookup.scala 11:37:@4199.4]
  assign _T_316 = _T_182 ? 2'h2 : 2'h0; // @[Lookup.scala 11:37:@4208.4]
  assign _T_317 = _T_178 ? 2'h0 : _T_316; // @[Lookup.scala 11:37:@4209.4]
  assign _T_318 = _T_174 ? 2'h0 : _T_317; // @[Lookup.scala 11:37:@4210.4]
  assign _T_319 = _T_170 ? 2'h0 : _T_318; // @[Lookup.scala 11:37:@4211.4]
  assign _T_320 = _T_166 ? 2'h2 : _T_319; // @[Lookup.scala 11:37:@4212.4]
  assign _T_321 = _T_162 ? 2'h2 : _T_320; // @[Lookup.scala 11:37:@4213.4]
  assign _T_322 = _T_158 ? 2'h0 : _T_321; // @[Lookup.scala 11:37:@4214.4]
  assign _T_323 = _T_154 ? 2'h0 : _T_322; // @[Lookup.scala 11:37:@4215.4]
  assign _T_324 = _T_150 ? 2'h0 : _T_323; // @[Lookup.scala 11:37:@4216.4]
  assign _T_325 = _T_146 ? 2'h0 : _T_324; // @[Lookup.scala 11:37:@4217.4]
  assign _T_326 = _T_142 ? 2'h0 : _T_325; // @[Lookup.scala 11:37:@4218.4]
  assign _T_327 = _T_138 ? 2'h0 : _T_326; // @[Lookup.scala 11:37:@4219.4]
  assign _T_328 = _T_134 ? 2'h0 : _T_327; // @[Lookup.scala 11:37:@4220.4]
  assign _T_329 = _T_130 ? 2'h0 : _T_328; // @[Lookup.scala 11:37:@4221.4]
  assign _T_330 = _T_126 ? 2'h0 : _T_329; // @[Lookup.scala 11:37:@4222.4]
  assign _T_331 = _T_122 ? 2'h0 : _T_330; // @[Lookup.scala 11:37:@4223.4]
  assign _T_332 = _T_118 ? 2'h0 : _T_331; // @[Lookup.scala 11:37:@4224.4]
  assign _T_333 = _T_114 ? 2'h0 : _T_332; // @[Lookup.scala 11:37:@4225.4]
  assign _T_334 = _T_110 ? 2'h0 : _T_333; // @[Lookup.scala 11:37:@4226.4]
  assign _T_335 = _T_106 ? 2'h0 : _T_334; // @[Lookup.scala 11:37:@4227.4]
  assign _T_336 = _T_102 ? 2'h0 : _T_335; // @[Lookup.scala 11:37:@4228.4]
  assign _T_337 = _T_98 ? 2'h0 : _T_336; // @[Lookup.scala 11:37:@4229.4]
  assign _T_338 = _T_94 ? 2'h0 : _T_337; // @[Lookup.scala 11:37:@4230.4]
  assign _T_339 = _T_90 ? 2'h0 : _T_338; // @[Lookup.scala 11:37:@4231.4]
  assign _T_340 = _T_86 ? 2'h0 : _T_339; // @[Lookup.scala 11:37:@4232.4]
  assign _T_341 = _T_82 ? 2'h0 : _T_340; // @[Lookup.scala 11:37:@4233.4]
  assign _T_342 = _T_78 ? 2'h0 : _T_341; // @[Lookup.scala 11:37:@4234.4]
  assign _T_343 = _T_74 ? 2'h0 : _T_342; // @[Lookup.scala 11:37:@4235.4]
  assign _T_344 = _T_70 ? 2'h0 : _T_343; // @[Lookup.scala 11:37:@4236.4]
  assign _T_345 = _T_66 ? 2'h0 : _T_344; // @[Lookup.scala 11:37:@4237.4]
  assign _T_346 = _T_62 ? 2'h0 : _T_345; // @[Lookup.scala 11:37:@4238.4]
  assign _T_347 = _T_58 ? 2'h0 : _T_346; // @[Lookup.scala 11:37:@4239.4]
  assign _T_348 = _T_54 ? 2'h0 : _T_347; // @[Lookup.scala 11:37:@4240.4]
  assign _T_349 = _T_50 ? 2'h0 : _T_348; // @[Lookup.scala 11:37:@4241.4]
  assign _T_350 = _T_46 ? 2'h1 : _T_349; // @[Lookup.scala 11:37:@4242.4]
  assign _T_351 = _T_42 ? 2'h0 : _T_350; // @[Lookup.scala 11:37:@4243.4]
  assign _T_352 = _T_38 ? 2'h0 : _T_351; // @[Lookup.scala 11:37:@4244.4]
  assign _T_353 = _T_34 ? 2'h0 : _T_352; // @[Lookup.scala 11:37:@4245.4]
  assign _T_354 = _T_30 ? 2'h0 : _T_353; // @[Lookup.scala 11:37:@4246.4]
  assign _T_355 = _T_26 ? 2'h0 : _T_354; // @[Lookup.scala 11:37:@4247.4]
  assign _T_356 = _T_22 ? 2'h0 : _T_355; // @[Lookup.scala 11:37:@4248.4]
  assign _T_357 = _T_18 ? 2'h0 : _T_356; // @[Lookup.scala 11:37:@4249.4]
  assign _T_371 = _T_158 ? 3'h3 : 3'h0; // @[Lookup.scala 11:37:@4264.4]
  assign _T_372 = _T_154 ? 3'h3 : _T_371; // @[Lookup.scala 11:37:@4265.4]
  assign _T_373 = _T_150 ? 3'h3 : _T_372; // @[Lookup.scala 11:37:@4266.4]
  assign _T_374 = _T_146 ? 3'h3 : _T_373; // @[Lookup.scala 11:37:@4267.4]
  assign _T_375 = _T_142 ? 3'h3 : _T_374; // @[Lookup.scala 11:37:@4268.4]
  assign _T_376 = _T_138 ? 3'h3 : _T_375; // @[Lookup.scala 11:37:@4269.4]
  assign _T_377 = _T_134 ? 3'h1 : _T_376; // @[Lookup.scala 11:37:@4270.4]
  assign _T_378 = _T_130 ? 3'h5 : _T_377; // @[Lookup.scala 11:37:@4271.4]
  assign _T_379 = _T_126 ? 3'h0 : _T_378; // @[Lookup.scala 11:37:@4272.4]
  assign _T_380 = _T_122 ? 3'h0 : _T_379; // @[Lookup.scala 11:37:@4273.4]
  assign _T_381 = _T_118 ? 3'h0 : _T_380; // @[Lookup.scala 11:37:@4274.4]
  assign _T_382 = _T_114 ? 3'h0 : _T_381; // @[Lookup.scala 11:37:@4275.4]
  assign _T_383 = _T_110 ? 3'h0 : _T_382; // @[Lookup.scala 11:37:@4276.4]
  assign _T_384 = _T_106 ? 3'h0 : _T_383; // @[Lookup.scala 11:37:@4277.4]
  assign _T_385 = _T_102 ? 3'h0 : _T_384; // @[Lookup.scala 11:37:@4278.4]
  assign _T_386 = _T_98 ? 3'h0 : _T_385; // @[Lookup.scala 11:37:@4279.4]
  assign _T_387 = _T_94 ? 3'h0 : _T_386; // @[Lookup.scala 11:37:@4280.4]
  assign _T_388 = _T_90 ? 3'h0 : _T_387; // @[Lookup.scala 11:37:@4281.4]
  assign _T_389 = _T_86 ? 3'h1 : _T_388; // @[Lookup.scala 11:37:@4282.4]
  assign _T_390 = _T_82 ? 3'h1 : _T_389; // @[Lookup.scala 11:37:@4283.4]
  assign _T_391 = _T_78 ? 3'h1 : _T_390; // @[Lookup.scala 11:37:@4284.4]
  assign _T_392 = _T_74 ? 3'h1 : _T_391; // @[Lookup.scala 11:37:@4285.4]
  assign _T_393 = _T_70 ? 3'h1 : _T_392; // @[Lookup.scala 11:37:@4286.4]
  assign _T_394 = _T_66 ? 3'h1 : _T_393; // @[Lookup.scala 11:37:@4287.4]
  assign _T_395 = _T_62 ? 3'h1 : _T_394; // @[Lookup.scala 11:37:@4288.4]
  assign _T_396 = _T_58 ? 3'h1 : _T_395; // @[Lookup.scala 11:37:@4289.4]
  assign _T_397 = _T_54 ? 3'h1 : _T_396; // @[Lookup.scala 11:37:@4290.4]
  assign _T_398 = _T_50 ? 3'h4 : _T_397; // @[Lookup.scala 11:37:@4291.4]
  assign _T_399 = _T_46 ? 3'h4 : _T_398; // @[Lookup.scala 11:37:@4292.4]
  assign _T_400 = _T_42 ? 3'h2 : _T_399; // @[Lookup.scala 11:37:@4293.4]
  assign _T_401 = _T_38 ? 3'h2 : _T_400; // @[Lookup.scala 11:37:@4294.4]
  assign _T_402 = _T_34 ? 3'h2 : _T_401; // @[Lookup.scala 11:37:@4295.4]
  assign _T_403 = _T_30 ? 3'h1 : _T_402; // @[Lookup.scala 11:37:@4296.4]
  assign _T_404 = _T_26 ? 3'h1 : _T_403; // @[Lookup.scala 11:37:@4297.4]
  assign _T_405 = _T_22 ? 3'h1 : _T_404; // @[Lookup.scala 11:37:@4298.4]
  assign _T_406 = _T_18 ? 3'h1 : _T_405; // @[Lookup.scala 11:37:@4299.4]
  assign _T_415 = _T_178 ? 1'h1 : _T_182; // @[Lookup.scala 11:37:@4309.4]
  assign _T_416 = _T_174 ? 1'h1 : _T_415; // @[Lookup.scala 11:37:@4310.4]
  assign _T_417 = _T_170 ? 1'h1 : _T_416; // @[Lookup.scala 11:37:@4311.4]
  assign _T_418 = _T_166 ? 1'h1 : _T_417; // @[Lookup.scala 11:37:@4312.4]
  assign _T_419 = _T_162 ? 1'h1 : _T_418; // @[Lookup.scala 11:37:@4313.4]
  assign _T_420 = _T_158 ? 1'h1 : _T_419; // @[Lookup.scala 11:37:@4314.4]
  assign _T_421 = _T_154 ? 1'h1 : _T_420; // @[Lookup.scala 11:37:@4315.4]
  assign _T_422 = _T_150 ? 1'h1 : _T_421; // @[Lookup.scala 11:37:@4316.4]
  assign _T_423 = _T_146 ? 1'h1 : _T_422; // @[Lookup.scala 11:37:@4317.4]
  assign _T_424 = _T_142 ? 1'h1 : _T_423; // @[Lookup.scala 11:37:@4318.4]
  assign _T_425 = _T_138 ? 1'h1 : _T_424; // @[Lookup.scala 11:37:@4319.4]
  assign _T_426 = _T_134 ? 1'h1 : _T_425; // @[Lookup.scala 11:37:@4320.4]
  assign _T_427 = _T_130 ? 1'h0 : _T_426; // @[Lookup.scala 11:37:@4321.4]
  assign _T_428 = _T_126 ? 1'h1 : _T_427; // @[Lookup.scala 11:37:@4322.4]
  assign _T_429 = _T_122 ? 1'h1 : _T_428; // @[Lookup.scala 11:37:@4323.4]
  assign _T_430 = _T_118 ? 1'h1 : _T_429; // @[Lookup.scala 11:37:@4324.4]
  assign _T_431 = _T_114 ? 1'h1 : _T_430; // @[Lookup.scala 11:37:@4325.4]
  assign _T_432 = _T_110 ? 1'h1 : _T_431; // @[Lookup.scala 11:37:@4326.4]
  assign _T_433 = _T_106 ? 1'h1 : _T_432; // @[Lookup.scala 11:37:@4327.4]
  assign _T_434 = _T_102 ? 1'h1 : _T_433; // @[Lookup.scala 11:37:@4328.4]
  assign _T_435 = _T_98 ? 1'h1 : _T_434; // @[Lookup.scala 11:37:@4329.4]
  assign _T_436 = _T_94 ? 1'h1 : _T_435; // @[Lookup.scala 11:37:@4330.4]
  assign _T_437 = _T_90 ? 1'h1 : _T_436; // @[Lookup.scala 11:37:@4331.4]
  assign _T_438 = _T_86 ? 1'h1 : _T_437; // @[Lookup.scala 11:37:@4332.4]
  assign _T_439 = _T_82 ? 1'h1 : _T_438; // @[Lookup.scala 11:37:@4333.4]
  assign _T_440 = _T_78 ? 1'h1 : _T_439; // @[Lookup.scala 11:37:@4334.4]
  assign _T_441 = _T_74 ? 1'h1 : _T_440; // @[Lookup.scala 11:37:@4335.4]
  assign _T_442 = _T_70 ? 1'h1 : _T_441; // @[Lookup.scala 11:37:@4336.4]
  assign _T_443 = _T_66 ? 1'h1 : _T_442; // @[Lookup.scala 11:37:@4337.4]
  assign _T_444 = _T_62 ? 1'h1 : _T_443; // @[Lookup.scala 11:37:@4338.4]
  assign _T_445 = _T_58 ? 1'h1 : _T_444; // @[Lookup.scala 11:37:@4339.4]
  assign _T_446 = _T_54 ? 1'h1 : _T_445; // @[Lookup.scala 11:37:@4340.4]
  assign _T_447 = _T_50 ? 1'h0 : _T_446; // @[Lookup.scala 11:37:@4341.4]
  assign _T_448 = _T_46 ? 1'h0 : _T_447; // @[Lookup.scala 11:37:@4342.4]
  assign _T_449 = _T_42 ? 1'h1 : _T_448; // @[Lookup.scala 11:37:@4343.4]
  assign _T_450 = _T_38 ? 1'h1 : _T_449; // @[Lookup.scala 11:37:@4344.4]
  assign _T_451 = _T_34 ? 1'h1 : _T_450; // @[Lookup.scala 11:37:@4345.4]
  assign _T_452 = _T_30 ? 1'h1 : _T_451; // @[Lookup.scala 11:37:@4346.4]
  assign _T_453 = _T_26 ? 1'h1 : _T_452; // @[Lookup.scala 11:37:@4347.4]
  assign _T_454 = _T_22 ? 1'h1 : _T_453; // @[Lookup.scala 11:37:@4348.4]
  assign _T_455 = _T_18 ? 1'h1 : _T_454; // @[Lookup.scala 11:37:@4349.4]
  assign _T_475 = _T_134 ? 1'h0 : _T_425; // @[Lookup.scala 11:37:@4370.4]
  assign _T_476 = _T_130 ? 1'h0 : _T_475; // @[Lookup.scala 11:37:@4371.4]
  assign _T_477 = _T_126 ? 1'h1 : _T_476; // @[Lookup.scala 11:37:@4372.4]
  assign _T_478 = _T_122 ? 1'h1 : _T_477; // @[Lookup.scala 11:37:@4373.4]
  assign _T_479 = _T_118 ? 1'h1 : _T_478; // @[Lookup.scala 11:37:@4374.4]
  assign _T_480 = _T_114 ? 1'h1 : _T_479; // @[Lookup.scala 11:37:@4375.4]
  assign _T_481 = _T_110 ? 1'h1 : _T_480; // @[Lookup.scala 11:37:@4376.4]
  assign _T_482 = _T_106 ? 1'h1 : _T_481; // @[Lookup.scala 11:37:@4377.4]
  assign _T_483 = _T_102 ? 1'h1 : _T_482; // @[Lookup.scala 11:37:@4378.4]
  assign _T_484 = _T_98 ? 1'h1 : _T_483; // @[Lookup.scala 11:37:@4379.4]
  assign _T_485 = _T_94 ? 1'h1 : _T_484; // @[Lookup.scala 11:37:@4380.4]
  assign _T_486 = _T_90 ? 1'h1 : _T_485; // @[Lookup.scala 11:37:@4381.4]
  assign _T_487 = _T_86 ? 1'h0 : _T_486; // @[Lookup.scala 11:37:@4382.4]
  assign _T_488 = _T_82 ? 1'h0 : _T_487; // @[Lookup.scala 11:37:@4383.4]
  assign _T_489 = _T_78 ? 1'h0 : _T_488; // @[Lookup.scala 11:37:@4384.4]
  assign _T_490 = _T_74 ? 1'h0 : _T_489; // @[Lookup.scala 11:37:@4385.4]
  assign _T_491 = _T_70 ? 1'h0 : _T_490; // @[Lookup.scala 11:37:@4386.4]
  assign _T_492 = _T_66 ? 1'h0 : _T_491; // @[Lookup.scala 11:37:@4387.4]
  assign _T_493 = _T_62 ? 1'h0 : _T_492; // @[Lookup.scala 11:37:@4388.4]
  assign _T_494 = _T_58 ? 1'h0 : _T_493; // @[Lookup.scala 11:37:@4389.4]
  assign _T_495 = _T_54 ? 1'h0 : _T_494; // @[Lookup.scala 11:37:@4390.4]
  assign _T_496 = _T_50 ? 1'h0 : _T_495; // @[Lookup.scala 11:37:@4391.4]
  assign _T_497 = _T_46 ? 1'h0 : _T_496; // @[Lookup.scala 11:37:@4392.4]
  assign _T_498 = _T_42 ? 1'h1 : _T_497; // @[Lookup.scala 11:37:@4393.4]
  assign _T_499 = _T_38 ? 1'h1 : _T_498; // @[Lookup.scala 11:37:@4394.4]
  assign _T_500 = _T_34 ? 1'h1 : _T_499; // @[Lookup.scala 11:37:@4395.4]
  assign _T_501 = _T_30 ? 1'h0 : _T_500; // @[Lookup.scala 11:37:@4396.4]
  assign _T_502 = _T_26 ? 1'h0 : _T_501; // @[Lookup.scala 11:37:@4397.4]
  assign _T_503 = _T_22 ? 1'h0 : _T_502; // @[Lookup.scala 11:37:@4398.4]
  assign _T_504 = _T_18 ? 1'h0 : _T_503; // @[Lookup.scala 11:37:@4399.4]
  assign _T_512 = _T_182 ? 4'ha : 4'h0; // @[Lookup.scala 11:37:@4408.4]
  assign _T_513 = _T_178 ? 4'ha : _T_512; // @[Lookup.scala 11:37:@4409.4]
  assign _T_514 = _T_174 ? 4'ha : _T_513; // @[Lookup.scala 11:37:@4410.4]
  assign _T_515 = _T_170 ? 4'ha : _T_514; // @[Lookup.scala 11:37:@4411.4]
  assign _T_516 = _T_166 ? 4'ha : _T_515; // @[Lookup.scala 11:37:@4412.4]
  assign _T_517 = _T_162 ? 4'ha : _T_516; // @[Lookup.scala 11:37:@4413.4]
  assign _T_518 = _T_158 ? 4'h0 : _T_517; // @[Lookup.scala 11:37:@4414.4]
  assign _T_519 = _T_154 ? 4'h0 : _T_518; // @[Lookup.scala 11:37:@4415.4]
  assign _T_520 = _T_150 ? 4'h0 : _T_519; // @[Lookup.scala 11:37:@4416.4]
  assign _T_521 = _T_146 ? 4'h0 : _T_520; // @[Lookup.scala 11:37:@4417.4]
  assign _T_522 = _T_142 ? 4'h0 : _T_521; // @[Lookup.scala 11:37:@4418.4]
  assign _T_523 = _T_138 ? 4'h0 : _T_522; // @[Lookup.scala 11:37:@4419.4]
  assign _T_524 = _T_134 ? 4'h0 : _T_523; // @[Lookup.scala 11:37:@4420.4]
  assign _T_525 = _T_130 ? 4'h0 : _T_524; // @[Lookup.scala 11:37:@4421.4]
  assign _T_526 = _T_126 ? 4'h3 : _T_525; // @[Lookup.scala 11:37:@4422.4]
  assign _T_527 = _T_122 ? 4'h4 : _T_526; // @[Lookup.scala 11:37:@4423.4]
  assign _T_528 = _T_118 ? 4'h7 : _T_527; // @[Lookup.scala 11:37:@4424.4]
  assign _T_529 = _T_114 ? 4'h6 : _T_528; // @[Lookup.scala 11:37:@4425.4]
  assign _T_530 = _T_110 ? 4'h5 : _T_529; // @[Lookup.scala 11:37:@4426.4]
  assign _T_531 = _T_106 ? 4'h9 : _T_530; // @[Lookup.scala 11:37:@4427.4]
  assign _T_532 = _T_102 ? 4'h8 : _T_531; // @[Lookup.scala 11:37:@4428.4]
  assign _T_533 = _T_98 ? 4'h1 : _T_532; // @[Lookup.scala 11:37:@4429.4]
  assign _T_534 = _T_94 ? 4'h0 : _T_533; // @[Lookup.scala 11:37:@4430.4]
  assign _T_535 = _T_90 ? 4'h2 : _T_534; // @[Lookup.scala 11:37:@4431.4]
  assign _T_536 = _T_86 ? 4'h3 : _T_535; // @[Lookup.scala 11:37:@4432.4]
  assign _T_537 = _T_82 ? 4'h4 : _T_536; // @[Lookup.scala 11:37:@4433.4]
  assign _T_538 = _T_78 ? 4'h2 : _T_537; // @[Lookup.scala 11:37:@4434.4]
  assign _T_539 = _T_74 ? 4'h9 : _T_538; // @[Lookup.scala 11:37:@4435.4]
  assign _T_540 = _T_70 ? 4'h8 : _T_539; // @[Lookup.scala 11:37:@4436.4]
  assign _T_541 = _T_66 ? 4'h7 : _T_540; // @[Lookup.scala 11:37:@4437.4]
  assign _T_542 = _T_62 ? 4'h6 : _T_541; // @[Lookup.scala 11:37:@4438.4]
  assign _T_543 = _T_58 ? 4'h5 : _T_542; // @[Lookup.scala 11:37:@4439.4]
  assign _T_544 = _T_54 ? 4'h0 : _T_543; // @[Lookup.scala 11:37:@4440.4]
  assign _T_545 = _T_50 ? 4'hb : _T_544; // @[Lookup.scala 11:37:@4441.4]
  assign _T_546 = _T_46 ? 4'h0 : _T_545; // @[Lookup.scala 11:37:@4442.4]
  assign _T_547 = _T_42 ? 4'h0 : _T_546; // @[Lookup.scala 11:37:@4443.4]
  assign _T_548 = _T_38 ? 4'h0 : _T_547; // @[Lookup.scala 11:37:@4444.4]
  assign _T_549 = _T_34 ? 4'h0 : _T_548; // @[Lookup.scala 11:37:@4445.4]
  assign _T_550 = _T_30 ? 4'h0 : _T_549; // @[Lookup.scala 11:37:@4446.4]
  assign _T_551 = _T_26 ? 4'h0 : _T_550; // @[Lookup.scala 11:37:@4447.4]
  assign _T_552 = _T_22 ? 4'h0 : _T_551; // @[Lookup.scala 11:37:@4448.4]
  assign _T_553 = _T_18 ? 4'h0 : _T_552; // @[Lookup.scala 11:37:@4449.4]
  assign _T_561 = _T_182 ? 2'h3 : 2'h0; // @[Lookup.scala 11:37:@4458.4]
  assign _T_562 = _T_178 ? 2'h3 : _T_561; // @[Lookup.scala 11:37:@4459.4]
  assign _T_563 = _T_174 ? 2'h3 : _T_562; // @[Lookup.scala 11:37:@4460.4]
  assign _T_564 = _T_170 ? 2'h3 : _T_563; // @[Lookup.scala 11:37:@4461.4]
  assign _T_565 = _T_166 ? 2'h3 : _T_564; // @[Lookup.scala 11:37:@4462.4]
  assign _T_566 = _T_162 ? 2'h3 : _T_565; // @[Lookup.scala 11:37:@4463.4]
  assign _T_567 = _T_158 ? 2'h0 : _T_566; // @[Lookup.scala 11:37:@4464.4]
  assign _T_568 = _T_154 ? 2'h0 : _T_567; // @[Lookup.scala 11:37:@4465.4]
  assign _T_569 = _T_150 ? 2'h0 : _T_568; // @[Lookup.scala 11:37:@4466.4]
  assign _T_570 = _T_146 ? 2'h0 : _T_569; // @[Lookup.scala 11:37:@4467.4]
  assign _T_571 = _T_142 ? 2'h0 : _T_570; // @[Lookup.scala 11:37:@4468.4]
  assign _T_572 = _T_138 ? 2'h0 : _T_571; // @[Lookup.scala 11:37:@4469.4]
  assign _T_573 = _T_134 ? 2'h2 : _T_572; // @[Lookup.scala 11:37:@4470.4]
  assign _T_574 = _T_130 ? 2'h2 : _T_573; // @[Lookup.scala 11:37:@4471.4]
  assign _T_575 = _T_126 ? 2'h0 : _T_574; // @[Lookup.scala 11:37:@4472.4]
  assign _T_576 = _T_122 ? 2'h0 : _T_575; // @[Lookup.scala 11:37:@4473.4]
  assign _T_577 = _T_118 ? 2'h0 : _T_576; // @[Lookup.scala 11:37:@4474.4]
  assign _T_578 = _T_114 ? 2'h0 : _T_577; // @[Lookup.scala 11:37:@4475.4]
  assign _T_579 = _T_110 ? 2'h0 : _T_578; // @[Lookup.scala 11:37:@4476.4]
  assign _T_580 = _T_106 ? 2'h0 : _T_579; // @[Lookup.scala 11:37:@4477.4]
  assign _T_581 = _T_102 ? 2'h0 : _T_580; // @[Lookup.scala 11:37:@4478.4]
  assign _T_582 = _T_98 ? 2'h0 : _T_581; // @[Lookup.scala 11:37:@4479.4]
  assign _T_583 = _T_94 ? 2'h0 : _T_582; // @[Lookup.scala 11:37:@4480.4]
  assign _T_584 = _T_90 ? 2'h0 : _T_583; // @[Lookup.scala 11:37:@4481.4]
  assign _T_585 = _T_86 ? 2'h0 : _T_584; // @[Lookup.scala 11:37:@4482.4]
  assign _T_586 = _T_82 ? 2'h0 : _T_585; // @[Lookup.scala 11:37:@4483.4]
  assign _T_587 = _T_78 ? 2'h0 : _T_586; // @[Lookup.scala 11:37:@4484.4]
  assign _T_588 = _T_74 ? 2'h0 : _T_587; // @[Lookup.scala 11:37:@4485.4]
  assign _T_589 = _T_70 ? 2'h0 : _T_588; // @[Lookup.scala 11:37:@4486.4]
  assign _T_590 = _T_66 ? 2'h0 : _T_589; // @[Lookup.scala 11:37:@4487.4]
  assign _T_591 = _T_62 ? 2'h0 : _T_590; // @[Lookup.scala 11:37:@4488.4]
  assign _T_592 = _T_58 ? 2'h0 : _T_591; // @[Lookup.scala 11:37:@4489.4]
  assign _T_593 = _T_54 ? 2'h0 : _T_592; // @[Lookup.scala 11:37:@4490.4]
  assign _T_594 = _T_50 ? 2'h0 : _T_593; // @[Lookup.scala 11:37:@4491.4]
  assign _T_595 = _T_46 ? 2'h0 : _T_594; // @[Lookup.scala 11:37:@4492.4]
  assign _T_596 = _T_42 ? 2'h0 : _T_595; // @[Lookup.scala 11:37:@4493.4]
  assign _T_597 = _T_38 ? 2'h0 : _T_596; // @[Lookup.scala 11:37:@4494.4]
  assign _T_598 = _T_34 ? 2'h0 : _T_597; // @[Lookup.scala 11:37:@4495.4]
  assign _T_599 = _T_30 ? 2'h1 : _T_598; // @[Lookup.scala 11:37:@4496.4]
  assign _T_600 = _T_26 ? 2'h1 : _T_599; // @[Lookup.scala 11:37:@4497.4]
  assign _T_601 = _T_22 ? 2'h1 : _T_600; // @[Lookup.scala 11:37:@4498.4]
  assign _T_602 = _T_18 ? 2'h1 : _T_601; // @[Lookup.scala 11:37:@4499.4]
  assign _T_616 = _T_158 ? 1'h0 : _T_419; // @[Lookup.scala 11:37:@4514.4]
  assign _T_617 = _T_154 ? 1'h0 : _T_616; // @[Lookup.scala 11:37:@4515.4]
  assign _T_618 = _T_150 ? 1'h0 : _T_617; // @[Lookup.scala 11:37:@4516.4]
  assign _T_619 = _T_146 ? 1'h0 : _T_618; // @[Lookup.scala 11:37:@4517.4]
  assign _T_620 = _T_142 ? 1'h0 : _T_619; // @[Lookup.scala 11:37:@4518.4]
  assign _T_621 = _T_138 ? 1'h0 : _T_620; // @[Lookup.scala 11:37:@4519.4]
  assign _T_622 = _T_134 ? 1'h1 : _T_621; // @[Lookup.scala 11:37:@4520.4]
  assign _T_623 = _T_130 ? 1'h1 : _T_622; // @[Lookup.scala 11:37:@4521.4]
  assign _T_624 = _T_126 ? 1'h1 : _T_623; // @[Lookup.scala 11:37:@4522.4]
  assign _T_625 = _T_122 ? 1'h1 : _T_624; // @[Lookup.scala 11:37:@4523.4]
  assign _T_626 = _T_118 ? 1'h1 : _T_625; // @[Lookup.scala 11:37:@4524.4]
  assign _T_627 = _T_114 ? 1'h1 : _T_626; // @[Lookup.scala 11:37:@4525.4]
  assign _T_628 = _T_110 ? 1'h1 : _T_627; // @[Lookup.scala 11:37:@4526.4]
  assign _T_629 = _T_106 ? 1'h1 : _T_628; // @[Lookup.scala 11:37:@4527.4]
  assign _T_630 = _T_102 ? 1'h1 : _T_629; // @[Lookup.scala 11:37:@4528.4]
  assign _T_631 = _T_98 ? 1'h1 : _T_630; // @[Lookup.scala 11:37:@4529.4]
  assign _T_632 = _T_94 ? 1'h1 : _T_631; // @[Lookup.scala 11:37:@4530.4]
  assign _T_633 = _T_90 ? 1'h1 : _T_632; // @[Lookup.scala 11:37:@4531.4]
  assign _T_634 = _T_86 ? 1'h1 : _T_633; // @[Lookup.scala 11:37:@4532.4]
  assign _T_635 = _T_82 ? 1'h1 : _T_634; // @[Lookup.scala 11:37:@4533.4]
  assign _T_636 = _T_78 ? 1'h1 : _T_635; // @[Lookup.scala 11:37:@4534.4]
  assign _T_637 = _T_74 ? 1'h1 : _T_636; // @[Lookup.scala 11:37:@4535.4]
  assign _T_638 = _T_70 ? 1'h1 : _T_637; // @[Lookup.scala 11:37:@4536.4]
  assign _T_639 = _T_66 ? 1'h1 : _T_638; // @[Lookup.scala 11:37:@4537.4]
  assign _T_640 = _T_62 ? 1'h1 : _T_639; // @[Lookup.scala 11:37:@4538.4]
  assign _T_641 = _T_58 ? 1'h1 : _T_640; // @[Lookup.scala 11:37:@4539.4]
  assign _T_642 = _T_54 ? 1'h1 : _T_641; // @[Lookup.scala 11:37:@4540.4]
  assign _T_643 = _T_50 ? 1'h1 : _T_642; // @[Lookup.scala 11:37:@4541.4]
  assign _T_644 = _T_46 ? 1'h1 : _T_643; // @[Lookup.scala 11:37:@4542.4]
  assign _T_645 = _T_42 ? 1'h0 : _T_644; // @[Lookup.scala 11:37:@4543.4]
  assign _T_646 = _T_38 ? 1'h0 : _T_645; // @[Lookup.scala 11:37:@4544.4]
  assign _T_647 = _T_34 ? 1'h0 : _T_646; // @[Lookup.scala 11:37:@4545.4]
  assign _T_648 = _T_30 ? 1'h1 : _T_647; // @[Lookup.scala 11:37:@4546.4]
  assign _T_649 = _T_26 ? 1'h1 : _T_648; // @[Lookup.scala 11:37:@4547.4]
  assign _T_650 = _T_22 ? 1'h1 : _T_649; // @[Lookup.scala 11:37:@4548.4]
  assign _T_651 = _T_18 ? 1'h1 : _T_650; // @[Lookup.scala 11:37:@4549.4]
  assign _T_653 = _T_206 ? 1'h0 : _T_210; // @[Lookup.scala 11:37:@4552.4]
  assign _T_654 = _T_202 ? 1'h0 : _T_653; // @[Lookup.scala 11:37:@4553.4]
  assign _T_655 = _T_198 ? 1'h0 : _T_654; // @[Lookup.scala 11:37:@4554.4]
  assign _T_656 = _T_194 ? 1'h0 : _T_655; // @[Lookup.scala 11:37:@4555.4]
  assign _T_657 = _T_190 ? 1'h0 : _T_656; // @[Lookup.scala 11:37:@4556.4]
  assign _T_658 = _T_186 ? 1'h0 : _T_657; // @[Lookup.scala 11:37:@4557.4]
  assign _T_659 = _T_182 ? 1'h0 : _T_658; // @[Lookup.scala 11:37:@4558.4]
  assign _T_660 = _T_178 ? 1'h0 : _T_659; // @[Lookup.scala 11:37:@4559.4]
  assign _T_661 = _T_174 ? 1'h0 : _T_660; // @[Lookup.scala 11:37:@4560.4]
  assign _T_662 = _T_170 ? 1'h0 : _T_661; // @[Lookup.scala 11:37:@4561.4]
  assign _T_663 = _T_166 ? 1'h0 : _T_662; // @[Lookup.scala 11:37:@4562.4]
  assign _T_664 = _T_162 ? 1'h0 : _T_663; // @[Lookup.scala 11:37:@4563.4]
  assign _T_665 = _T_158 ? 1'h0 : _T_664; // @[Lookup.scala 11:37:@4564.4]
  assign _T_666 = _T_154 ? 1'h0 : _T_665; // @[Lookup.scala 11:37:@4565.4]
  assign _T_667 = _T_150 ? 1'h0 : _T_666; // @[Lookup.scala 11:37:@4566.4]
  assign _T_668 = _T_146 ? 1'h0 : _T_667; // @[Lookup.scala 11:37:@4567.4]
  assign _T_669 = _T_142 ? 1'h0 : _T_668; // @[Lookup.scala 11:37:@4568.4]
  assign _T_670 = _T_138 ? 1'h0 : _T_669; // @[Lookup.scala 11:37:@4569.4]
  assign _T_671 = _T_134 ? 1'h0 : _T_670; // @[Lookup.scala 11:37:@4570.4]
  assign _T_672 = _T_130 ? 1'h0 : _T_671; // @[Lookup.scala 11:37:@4571.4]
  assign _T_673 = _T_126 ? 1'h0 : _T_672; // @[Lookup.scala 11:37:@4572.4]
  assign _T_674 = _T_122 ? 1'h0 : _T_673; // @[Lookup.scala 11:37:@4573.4]
  assign _T_675 = _T_118 ? 1'h0 : _T_674; // @[Lookup.scala 11:37:@4574.4]
  assign _T_676 = _T_114 ? 1'h0 : _T_675; // @[Lookup.scala 11:37:@4575.4]
  assign _T_677 = _T_110 ? 1'h0 : _T_676; // @[Lookup.scala 11:37:@4576.4]
  assign _T_678 = _T_106 ? 1'h0 : _T_677; // @[Lookup.scala 11:37:@4577.4]
  assign _T_679 = _T_102 ? 1'h0 : _T_678; // @[Lookup.scala 11:37:@4578.4]
  assign _T_680 = _T_98 ? 1'h0 : _T_679; // @[Lookup.scala 11:37:@4579.4]
  assign _T_681 = _T_94 ? 1'h0 : _T_680; // @[Lookup.scala 11:37:@4580.4]
  assign _T_682 = _T_90 ? 1'h0 : _T_681; // @[Lookup.scala 11:37:@4581.4]
  assign _T_683 = _T_86 ? 1'h0 : _T_682; // @[Lookup.scala 11:37:@4582.4]
  assign _T_684 = _T_82 ? 1'h0 : _T_683; // @[Lookup.scala 11:37:@4583.4]
  assign _T_685 = _T_78 ? 1'h0 : _T_684; // @[Lookup.scala 11:37:@4584.4]
  assign _T_686 = _T_74 ? 1'h0 : _T_685; // @[Lookup.scala 11:37:@4585.4]
  assign _T_687 = _T_70 ? 1'h0 : _T_686; // @[Lookup.scala 11:37:@4586.4]
  assign _T_688 = _T_66 ? 1'h0 : _T_687; // @[Lookup.scala 11:37:@4587.4]
  assign _T_689 = _T_62 ? 1'h0 : _T_688; // @[Lookup.scala 11:37:@4588.4]
  assign _T_690 = _T_58 ? 1'h0 : _T_689; // @[Lookup.scala 11:37:@4589.4]
  assign _T_691 = _T_54 ? 1'h0 : _T_690; // @[Lookup.scala 11:37:@4590.4]
  assign _T_692 = _T_50 ? 1'h0 : _T_691; // @[Lookup.scala 11:37:@4591.4]
  assign _T_693 = _T_46 ? 1'h0 : _T_692; // @[Lookup.scala 11:37:@4592.4]
  assign _T_694 = _T_42 ? 1'h1 : _T_693; // @[Lookup.scala 11:37:@4593.4]
  assign _T_695 = _T_38 ? 1'h1 : _T_694; // @[Lookup.scala 11:37:@4594.4]
  assign _T_696 = _T_34 ? 1'h1 : _T_695; // @[Lookup.scala 11:37:@4595.4]
  assign _T_697 = _T_30 ? 1'h1 : _T_696; // @[Lookup.scala 11:37:@4596.4]
  assign _T_698 = _T_26 ? 1'h1 : _T_697; // @[Lookup.scala 11:37:@4597.4]
  assign _T_699 = _T_22 ? 1'h1 : _T_698; // @[Lookup.scala 11:37:@4598.4]
  assign _T_700 = _T_18 ? 1'h1 : _T_699; // @[Lookup.scala 11:37:@4599.4]
  assign _T_744 = _T_38 ? 1'h1 : _T_42; // @[Lookup.scala 11:37:@4644.4]
  assign _T_745 = _T_34 ? 1'h1 : _T_744; // @[Lookup.scala 11:37:@4645.4]
  assign _T_746 = _T_30 ? 1'h0 : _T_745; // @[Lookup.scala 11:37:@4646.4]
  assign _T_747 = _T_26 ? 1'h0 : _T_746; // @[Lookup.scala 11:37:@4647.4]
  assign _T_748 = _T_22 ? 1'h0 : _T_747; // @[Lookup.scala 11:37:@4648.4]
  assign _T_749 = _T_18 ? 1'h0 : _T_748; // @[Lookup.scala 11:37:@4649.4]
  assign _T_792 = _T_42 ? 3'h2 : 3'h0; // @[Lookup.scala 11:37:@4693.4]
  assign _T_793 = _T_38 ? 3'h1 : _T_792; // @[Lookup.scala 11:37:@4694.4]
  assign _T_794 = _T_34 ? 3'h3 : _T_793; // @[Lookup.scala 11:37:@4695.4]
  assign _T_795 = _T_30 ? 3'h6 : _T_794; // @[Lookup.scala 11:37:@4696.4]
  assign _T_796 = _T_26 ? 3'h2 : _T_795; // @[Lookup.scala 11:37:@4697.4]
  assign _T_797 = _T_22 ? 3'h5 : _T_796; // @[Lookup.scala 11:37:@4698.4]
  assign _T_798 = _T_18 ? 3'h1 : _T_797; // @[Lookup.scala 11:37:@4699.4]
  assign _T_802 = _T_198 ? 3'h4 : 3'h0; // @[Lookup.scala 11:37:@4704.4]
  assign _T_803 = _T_194 ? 3'h4 : _T_802; // @[Lookup.scala 11:37:@4705.4]
  assign _T_804 = _T_190 ? 3'h4 : _T_803; // @[Lookup.scala 11:37:@4706.4]
  assign _T_805 = _T_186 ? 3'h4 : _T_804; // @[Lookup.scala 11:37:@4707.4]
  assign _T_806 = _T_182 ? 3'h3 : _T_805; // @[Lookup.scala 11:37:@4708.4]
  assign _T_807 = _T_178 ? 3'h3 : _T_806; // @[Lookup.scala 11:37:@4709.4]
  assign _T_808 = _T_174 ? 3'h2 : _T_807; // @[Lookup.scala 11:37:@4710.4]
  assign _T_809 = _T_170 ? 3'h1 : _T_808; // @[Lookup.scala 11:37:@4711.4]
  assign _T_810 = _T_166 ? 3'h2 : _T_809; // @[Lookup.scala 11:37:@4712.4]
  assign _T_811 = _T_162 ? 3'h1 : _T_810; // @[Lookup.scala 11:37:@4713.4]
  assign _T_812 = _T_158 ? 3'h0 : _T_811; // @[Lookup.scala 11:37:@4714.4]
  assign _T_813 = _T_154 ? 3'h0 : _T_812; // @[Lookup.scala 11:37:@4715.4]
  assign _T_814 = _T_150 ? 3'h0 : _T_813; // @[Lookup.scala 11:37:@4716.4]
  assign _T_815 = _T_146 ? 3'h0 : _T_814; // @[Lookup.scala 11:37:@4717.4]
  assign _T_816 = _T_142 ? 3'h0 : _T_815; // @[Lookup.scala 11:37:@4718.4]
  assign _T_817 = _T_138 ? 3'h0 : _T_816; // @[Lookup.scala 11:37:@4719.4]
  assign _T_818 = _T_134 ? 3'h0 : _T_817; // @[Lookup.scala 11:37:@4720.4]
  assign _T_819 = _T_130 ? 3'h0 : _T_818; // @[Lookup.scala 11:37:@4721.4]
  assign _T_820 = _T_126 ? 3'h0 : _T_819; // @[Lookup.scala 11:37:@4722.4]
  assign _T_821 = _T_122 ? 3'h0 : _T_820; // @[Lookup.scala 11:37:@4723.4]
  assign _T_822 = _T_118 ? 3'h0 : _T_821; // @[Lookup.scala 11:37:@4724.4]
  assign _T_823 = _T_114 ? 3'h0 : _T_822; // @[Lookup.scala 11:37:@4725.4]
  assign _T_824 = _T_110 ? 3'h0 : _T_823; // @[Lookup.scala 11:37:@4726.4]
  assign _T_825 = _T_106 ? 3'h0 : _T_824; // @[Lookup.scala 11:37:@4727.4]
  assign _T_826 = _T_102 ? 3'h0 : _T_825; // @[Lookup.scala 11:37:@4728.4]
  assign _T_827 = _T_98 ? 3'h0 : _T_826; // @[Lookup.scala 11:37:@4729.4]
  assign _T_828 = _T_94 ? 3'h0 : _T_827; // @[Lookup.scala 11:37:@4730.4]
  assign _T_829 = _T_90 ? 3'h0 : _T_828; // @[Lookup.scala 11:37:@4731.4]
  assign _T_830 = _T_86 ? 3'h0 : _T_829; // @[Lookup.scala 11:37:@4732.4]
  assign _T_831 = _T_82 ? 3'h0 : _T_830; // @[Lookup.scala 11:37:@4733.4]
  assign _T_832 = _T_78 ? 3'h0 : _T_831; // @[Lookup.scala 11:37:@4734.4]
  assign _T_833 = _T_74 ? 3'h0 : _T_832; // @[Lookup.scala 11:37:@4735.4]
  assign _T_834 = _T_70 ? 3'h0 : _T_833; // @[Lookup.scala 11:37:@4736.4]
  assign _T_835 = _T_66 ? 3'h0 : _T_834; // @[Lookup.scala 11:37:@4737.4]
  assign _T_836 = _T_62 ? 3'h0 : _T_835; // @[Lookup.scala 11:37:@4738.4]
  assign _T_837 = _T_58 ? 3'h0 : _T_836; // @[Lookup.scala 11:37:@4739.4]
  assign _T_838 = _T_54 ? 3'h0 : _T_837; // @[Lookup.scala 11:37:@4740.4]
  assign _T_839 = _T_50 ? 3'h0 : _T_838; // @[Lookup.scala 11:37:@4741.4]
  assign _T_840 = _T_46 ? 3'h0 : _T_839; // @[Lookup.scala 11:37:@4742.4]
  assign _T_841 = _T_42 ? 3'h0 : _T_840; // @[Lookup.scala 11:37:@4743.4]
  assign _T_842 = _T_38 ? 3'h0 : _T_841; // @[Lookup.scala 11:37:@4744.4]
  assign _T_843 = _T_34 ? 3'h0 : _T_842; // @[Lookup.scala 11:37:@4745.4]
  assign _T_844 = _T_30 ? 3'h0 : _T_843; // @[Lookup.scala 11:37:@4746.4]
  assign _T_845 = _T_26 ? 3'h0 : _T_844; // @[Lookup.scala 11:37:@4747.4]
  assign _T_846 = _T_22 ? 3'h0 : _T_845; // @[Lookup.scala 11:37:@4748.4]
  assign _T_847 = _T_18 ? 3'h0 : _T_846; // @[Lookup.scala 11:37:@4749.4]
  assign _T_850 = _T_202 ? 1'h0 : _T_206; // @[Lookup.scala 11:37:@4753.4]
  assign _T_851 = _T_198 ? 1'h0 : _T_850; // @[Lookup.scala 11:37:@4754.4]
  assign _T_852 = _T_194 ? 1'h0 : _T_851; // @[Lookup.scala 11:37:@4755.4]
  assign _T_853 = _T_190 ? 1'h0 : _T_852; // @[Lookup.scala 11:37:@4756.4]
  assign _T_854 = _T_186 ? 1'h0 : _T_853; // @[Lookup.scala 11:37:@4757.4]
  assign _T_855 = _T_182 ? 1'h0 : _T_854; // @[Lookup.scala 11:37:@4758.4]
  assign _T_856 = _T_178 ? 1'h0 : _T_855; // @[Lookup.scala 11:37:@4759.4]
  assign _T_857 = _T_174 ? 1'h0 : _T_856; // @[Lookup.scala 11:37:@4760.4]
  assign _T_858 = _T_170 ? 1'h0 : _T_857; // @[Lookup.scala 11:37:@4761.4]
  assign _T_859 = _T_166 ? 1'h0 : _T_858; // @[Lookup.scala 11:37:@4762.4]
  assign _T_860 = _T_162 ? 1'h0 : _T_859; // @[Lookup.scala 11:37:@4763.4]
  assign _T_861 = _T_158 ? 1'h0 : _T_860; // @[Lookup.scala 11:37:@4764.4]
  assign _T_862 = _T_154 ? 1'h0 : _T_861; // @[Lookup.scala 11:37:@4765.4]
  assign _T_863 = _T_150 ? 1'h0 : _T_862; // @[Lookup.scala 11:37:@4766.4]
  assign _T_864 = _T_146 ? 1'h0 : _T_863; // @[Lookup.scala 11:37:@4767.4]
  assign _T_865 = _T_142 ? 1'h0 : _T_864; // @[Lookup.scala 11:37:@4768.4]
  assign _T_866 = _T_138 ? 1'h0 : _T_865; // @[Lookup.scala 11:37:@4769.4]
  assign _T_867 = _T_134 ? 1'h0 : _T_866; // @[Lookup.scala 11:37:@4770.4]
  assign _T_868 = _T_130 ? 1'h0 : _T_867; // @[Lookup.scala 11:37:@4771.4]
  assign _T_869 = _T_126 ? 1'h0 : _T_868; // @[Lookup.scala 11:37:@4772.4]
  assign _T_870 = _T_122 ? 1'h0 : _T_869; // @[Lookup.scala 11:37:@4773.4]
  assign _T_871 = _T_118 ? 1'h0 : _T_870; // @[Lookup.scala 11:37:@4774.4]
  assign _T_872 = _T_114 ? 1'h0 : _T_871; // @[Lookup.scala 11:37:@4775.4]
  assign _T_873 = _T_110 ? 1'h0 : _T_872; // @[Lookup.scala 11:37:@4776.4]
  assign _T_874 = _T_106 ? 1'h0 : _T_873; // @[Lookup.scala 11:37:@4777.4]
  assign _T_875 = _T_102 ? 1'h0 : _T_874; // @[Lookup.scala 11:37:@4778.4]
  assign _T_876 = _T_98 ? 1'h0 : _T_875; // @[Lookup.scala 11:37:@4779.4]
  assign _T_877 = _T_94 ? 1'h0 : _T_876; // @[Lookup.scala 11:37:@4780.4]
  assign _T_878 = _T_90 ? 1'h0 : _T_877; // @[Lookup.scala 11:37:@4781.4]
  assign _T_879 = _T_86 ? 1'h0 : _T_878; // @[Lookup.scala 11:37:@4782.4]
  assign _T_880 = _T_82 ? 1'h0 : _T_879; // @[Lookup.scala 11:37:@4783.4]
  assign _T_881 = _T_78 ? 1'h0 : _T_880; // @[Lookup.scala 11:37:@4784.4]
  assign _T_882 = _T_74 ? 1'h0 : _T_881; // @[Lookup.scala 11:37:@4785.4]
  assign _T_883 = _T_70 ? 1'h0 : _T_882; // @[Lookup.scala 11:37:@4786.4]
  assign _T_884 = _T_66 ? 1'h0 : _T_883; // @[Lookup.scala 11:37:@4787.4]
  assign _T_885 = _T_62 ? 1'h0 : _T_884; // @[Lookup.scala 11:37:@4788.4]
  assign _T_886 = _T_58 ? 1'h0 : _T_885; // @[Lookup.scala 11:37:@4789.4]
  assign _T_887 = _T_54 ? 1'h0 : _T_886; // @[Lookup.scala 11:37:@4790.4]
  assign _T_888 = _T_50 ? 1'h0 : _T_887; // @[Lookup.scala 11:37:@4791.4]
  assign _T_889 = _T_46 ? 1'h0 : _T_888; // @[Lookup.scala 11:37:@4792.4]
  assign _T_890 = _T_42 ? 1'h0 : _T_889; // @[Lookup.scala 11:37:@4793.4]
  assign _T_891 = _T_38 ? 1'h0 : _T_890; // @[Lookup.scala 11:37:@4794.4]
  assign _T_892 = _T_34 ? 1'h0 : _T_891; // @[Lookup.scala 11:37:@4795.4]
  assign _T_893 = _T_30 ? 1'h0 : _T_892; // @[Lookup.scala 11:37:@4796.4]
  assign _T_894 = _T_26 ? 1'h0 : _T_893; // @[Lookup.scala 11:37:@4797.4]
  assign _T_895 = _T_22 ? 1'h0 : _T_894; // @[Lookup.scala 11:37:@4798.4]
  assign _T_896 = _T_18 ? 1'h0 : _T_895; // @[Lookup.scala 11:37:@4799.4]
  assign _T_899 = io_inst[19:15]; // @[InstDecoder.scala 130:31:@4816.4]
  assign _T_901 = io_inst[11:7]; // @[InstDecoder.scala 132:31:@4820.4]
  assign func = io_inst[6:2]; // @[InstDecoder.scala 134:21:@4822.4]
  assign _T_905 = func == 5'h1b; // @[InstDecoder.scala 136:38:@4825.4]
  assign _T_907 = func == 5'h19; // @[InstDecoder.scala 137:39:@4826.4]
  assign _T_908 = _T_905 | _T_907; // @[InstDecoder.scala 141:32:@4827.4]
  assign _T_910 = io_cinfo_wbaddr == 5'h1; // @[InstDecoder.scala 135:37:@4828.4]
  assign _T_912 = io_cinfo_wbaddr == 5'h5; // @[InstDecoder.scala 135:53:@4829.4]
  assign _T_913 = _T_910 | _T_912; // @[InstDecoder.scala 135:45:@4830.4]
  assign _GEN_0 = {{4'd0}, _T_907}; // @[InstDecoder.scala 142:24:@4834.4]
  assign _T_917 = func == _GEN_0; // @[InstDecoder.scala 142:24:@4834.4]
  assign _T_919 = io_cinfo_rs1_addr == 5'h1; // @[InstDecoder.scala 135:37:@4835.4]
  assign _T_921 = io_cinfo_rs1_addr == 5'h5; // @[InstDecoder.scala 135:53:@4836.4]
  assign _T_922 = _T_919 | _T_921; // @[InstDecoder.scala 135:45:@4837.4]
  assign _T_923 = _T_917 & _T_922; // @[InstDecoder.scala 142:41:@4838.4]
  assign _T_930 = _T_913 == 1'h0; // @[InstDecoder.scala 143:6:@4842.4]
  assign _T_931 = io_cinfo_rs1_addr != io_cinfo_wbaddr; // @[InstDecoder.scala 143:50:@4843.4]
  assign _T_932 = _T_930 | _T_931; // @[InstDecoder.scala 143:29:@4844.4]
  assign imm_itype = io_inst[31:20]; // @[InstDecoder.scala 146:27:@4847.4]
  assign _T_934 = io_inst[31:25]; // @[InstDecoder.scala 147:31:@4848.4]
  assign imm_stype = {_T_934,_T_901}; // @[Cat.scala 30:58:@4850.4]
  assign _T_936 = io_inst[31]; // @[InstDecoder.scala 148:31:@4851.4]
  assign _T_937 = io_inst[7]; // @[InstDecoder.scala 148:44:@4852.4]
  assign _T_938 = io_inst[30:25]; // @[InstDecoder.scala 148:56:@4853.4]
  assign _T_939 = io_inst[11:8]; // @[InstDecoder.scala 148:73:@4854.4]
  assign imm_sbtype = {_T_936,_T_937,_T_938,_T_939}; // @[Cat.scala 30:58:@4857.4]
  assign imm_utype = io_inst[31:12]; // @[InstDecoder.scala 149:27:@4858.4]
  assign _T_943 = io_inst[19:12]; // @[InstDecoder.scala 150:44:@4860.4]
  assign _T_944 = io_inst[20]; // @[InstDecoder.scala 150:60:@4861.4]
  assign _T_945 = io_inst[30:21]; // @[InstDecoder.scala 150:73:@4862.4]
  assign imm_ujtype = {_T_936,_T_943,_T_944,_T_945}; // @[Cat.scala 30:58:@4865.4]
  assign _T_948 = imm_itype[11]; // @[InstDecoder.scala 153:43:@4866.4]
  assign _T_952 = _T_948 ? 20'hfffff : 20'h0; // @[Bitwise.scala 72:12:@4868.4]
  assign _T_954 = imm_stype[11]; // @[InstDecoder.scala 154:43:@4871.4]
  assign _T_958 = _T_954 ? 20'hfffff : 20'h0; // @[Bitwise.scala 72:12:@4873.4]
  assign _T_960 = imm_sbtype[11]; // @[InstDecoder.scala 155:44:@4876.4]
  assign _T_964 = _T_960 ? 19'h7ffff : 19'h0; // @[Bitwise.scala 72:12:@4878.4]
  assign _T_966 = {_T_964,_T_936,_T_937,_T_938,_T_939}; // @[Cat.scala 30:58:@4879.4]
  assign _T_974 = imm_ujtype[19]; // @[InstDecoder.scala 157:44:@4885.4]
  assign _T_978 = _T_974 ? 11'h7ff : 11'h0; // @[Bitwise.scala 72:12:@4887.4]
  assign _T_980 = {_T_978,_T_936,_T_943,_T_944,_T_945}; // @[Cat.scala 30:58:@4888.4]
  assign io_cinfo_br_type = _T_14 ? 4'h0 : _T_308; // @[InstDecoder.scala 115:20:@4801.4]
  assign io_cinfo_op1_sel = _T_14 ? 2'h0 : _T_357; // @[InstDecoder.scala 116:20:@4802.4]
  assign io_cinfo_op2_sel = _T_14 ? 3'h1 : _T_406; // @[InstDecoder.scala 117:20:@4803.4]
  assign io_cinfo_rs1_oen = _T_14 ? 1'h1 : _T_455; // @[InstDecoder.scala 118:20:@4804.4]
  assign io_cinfo_rs2_oen = _T_14 ? 1'h0 : _T_504; // @[InstDecoder.scala 119:20:@4805.4]
  assign io_cinfo_alu_fun = _T_14 ? 4'h0 : _T_553; // @[InstDecoder.scala 120:20:@4806.4]
  assign io_cinfo_wb_sel = _T_14 ? 2'h1 : _T_602; // @[InstDecoder.scala 121:20:@4807.4]
  assign io_cinfo_rf_wen = _T_14 ? 1'h1 : _T_651; // @[InstDecoder.scala 122:20:@4808.4]
  assign io_cinfo_mem_en = _T_14 ? 1'h1 : _T_700; // @[InstDecoder.scala 123:20:@4809.4]
  assign io_cinfo_mem_fcn = _T_14 ? 1'h0 : _T_749; // @[InstDecoder.scala 124:20:@4810.4]
  assign io_cinfo_mem_typ = _T_14 ? 3'h3 : _T_798; // @[InstDecoder.scala 125:20:@4811.4]
  assign io_cinfo_csr_cmd = _T_14 ? 3'h0 : _T_847; // @[InstDecoder.scala 126:20:@4812.4]
  assign io_cinfo_illegal = signals_0 == 1'h0; // @[InstDecoder.scala 127:20:@4814.4]
  assign io_cinfo_fencei = _T_14 ? 1'h0 : _T_896; // @[InstDecoder.scala 128:20:@4815.4]
  assign io_cinfo_is_branch = func == 5'h18; // @[InstDecoder.scala 139:22:@4824.4]
  assign io_cinfo_push = _T_908 & _T_913; // @[InstDecoder.scala 141:17:@4832.4]
  assign io_cinfo_pop = _T_923 & _T_932; // @[InstDecoder.scala 142:16:@4846.4]
  assign io_cinfo_rs1_addr = io_inst[19:15]; // @[InstDecoder.scala 130:21:@4817.4]
  assign io_cinfo_rs2_addr = io_inst[24:20]; // @[InstDecoder.scala 131:21:@4819.4]
  assign io_cinfo_wbaddr = io_inst[11:7]; // @[InstDecoder.scala 132:21:@4821.4]
  assign io_dinfo_imm_i = {_T_952,imm_itype}; // @[InstDecoder.scala 153:19:@4870.4]
  assign io_dinfo_imm_s = {_T_958,imm_stype}; // @[InstDecoder.scala 154:19:@4875.4]
  assign io_dinfo_imm_sb = {_T_966,1'h0}; // @[InstDecoder.scala 155:19:@4881.4]
  assign io_dinfo_imm_u = {imm_utype,12'h0}; // @[InstDecoder.scala 156:19:@4884.4]
  assign io_dinfo_imm_uj = {_T_980,1'h0}; // @[InstDecoder.scala 157:19:@4890.4]
  assign io_dinfo_imm_z = {27'h0,_T_899}; // @[InstDecoder.scala 158:19:@4894.4]
endmodule